magic
tech sky130A
magscale 1 2
timestamp 1647795232
<< obsli1 >>
rect 949 1581 253707 304657
<< obsm1 >>
rect 198 1096 254274 304688
<< metal2 >>
rect 1122 306339 1178 307139
rect 3330 306339 3386 307139
rect 5538 306339 5594 307139
rect 7746 306339 7802 307139
rect 10046 306339 10102 307139
rect 12254 306339 12310 307139
rect 14462 306339 14518 307139
rect 16670 306339 16726 307139
rect 18970 306339 19026 307139
rect 21178 306339 21234 307139
rect 23386 306339 23442 307139
rect 25594 306339 25650 307139
rect 27894 306339 27950 307139
rect 30102 306339 30158 307139
rect 32310 306339 32366 307139
rect 34610 306339 34666 307139
rect 36818 306339 36874 307139
rect 39026 306339 39082 307139
rect 41234 306339 41290 307139
rect 43534 306339 43590 307139
rect 45742 306339 45798 307139
rect 47950 306339 48006 307139
rect 50158 306339 50214 307139
rect 52458 306339 52514 307139
rect 54666 306339 54722 307139
rect 56874 306339 56930 307139
rect 59174 306339 59230 307139
rect 61382 306339 61438 307139
rect 63590 306339 63646 307139
rect 65798 306339 65854 307139
rect 68098 306339 68154 307139
rect 70306 306339 70362 307139
rect 72514 306339 72570 307139
rect 74722 306339 74778 307139
rect 77022 306339 77078 307139
rect 79230 306339 79286 307139
rect 81438 306339 81494 307139
rect 83738 306339 83794 307139
rect 85946 306339 86002 307139
rect 88154 306339 88210 307139
rect 90362 306339 90418 307139
rect 92662 306339 92718 307139
rect 94870 306339 94926 307139
rect 97078 306339 97134 307139
rect 99286 306339 99342 307139
rect 101586 306339 101642 307139
rect 103794 306339 103850 307139
rect 106002 306339 106058 307139
rect 108302 306339 108358 307139
rect 110510 306339 110566 307139
rect 112718 306339 112774 307139
rect 114926 306339 114982 307139
rect 117226 306339 117282 307139
rect 119434 306339 119490 307139
rect 121642 306339 121698 307139
rect 123850 306339 123906 307139
rect 126150 306339 126206 307139
rect 128358 306339 128414 307139
rect 130566 306339 130622 307139
rect 132866 306339 132922 307139
rect 135074 306339 135130 307139
rect 137282 306339 137338 307139
rect 139490 306339 139546 307139
rect 141790 306339 141846 307139
rect 143998 306339 144054 307139
rect 146206 306339 146262 307139
rect 148414 306339 148470 307139
rect 150714 306339 150770 307139
rect 152922 306339 152978 307139
rect 155130 306339 155186 307139
rect 157430 306339 157486 307139
rect 159638 306339 159694 307139
rect 161846 306339 161902 307139
rect 164054 306339 164110 307139
rect 166354 306339 166410 307139
rect 168562 306339 168618 307139
rect 170770 306339 170826 307139
rect 172978 306339 173034 307139
rect 175278 306339 175334 307139
rect 177486 306339 177542 307139
rect 179694 306339 179750 307139
rect 181994 306339 182050 307139
rect 184202 306339 184258 307139
rect 186410 306339 186466 307139
rect 188618 306339 188674 307139
rect 190918 306339 190974 307139
rect 193126 306339 193182 307139
rect 195334 306339 195390 307139
rect 197542 306339 197598 307139
rect 199842 306339 199898 307139
rect 202050 306339 202106 307139
rect 204258 306339 204314 307139
rect 206558 306339 206614 307139
rect 208766 306339 208822 307139
rect 210974 306339 211030 307139
rect 213182 306339 213238 307139
rect 215482 306339 215538 307139
rect 217690 306339 217746 307139
rect 219898 306339 219954 307139
rect 222106 306339 222162 307139
rect 224406 306339 224462 307139
rect 226614 306339 226670 307139
rect 228822 306339 228878 307139
rect 231122 306339 231178 307139
rect 233330 306339 233386 307139
rect 235538 306339 235594 307139
rect 237746 306339 237802 307139
rect 240046 306339 240102 307139
rect 242254 306339 242310 307139
rect 244462 306339 244518 307139
rect 246670 306339 246726 307139
rect 248970 306339 249026 307139
rect 251178 306339 251234 307139
rect 253386 306339 253442 307139
rect 202 0 258 800
rect 662 0 718 800
rect 1214 0 1270 800
rect 1674 0 1730 800
rect 2226 0 2282 800
rect 2778 0 2834 800
rect 3238 0 3294 800
rect 3790 0 3846 800
rect 4250 0 4306 800
rect 4802 0 4858 800
rect 5354 0 5410 800
rect 5814 0 5870 800
rect 6366 0 6422 800
rect 6826 0 6882 800
rect 7378 0 7434 800
rect 7930 0 7986 800
rect 8390 0 8446 800
rect 8942 0 8998 800
rect 9494 0 9550 800
rect 9954 0 10010 800
rect 10506 0 10562 800
rect 10966 0 11022 800
rect 11518 0 11574 800
rect 12070 0 12126 800
rect 12530 0 12586 800
rect 13082 0 13138 800
rect 13542 0 13598 800
rect 14094 0 14150 800
rect 14646 0 14702 800
rect 15106 0 15162 800
rect 15658 0 15714 800
rect 16118 0 16174 800
rect 16670 0 16726 800
rect 17222 0 17278 800
rect 17682 0 17738 800
rect 18234 0 18290 800
rect 18786 0 18842 800
rect 19246 0 19302 800
rect 19798 0 19854 800
rect 20258 0 20314 800
rect 20810 0 20866 800
rect 21362 0 21418 800
rect 21822 0 21878 800
rect 22374 0 22430 800
rect 22834 0 22890 800
rect 23386 0 23442 800
rect 23938 0 23994 800
rect 24398 0 24454 800
rect 24950 0 25006 800
rect 25502 0 25558 800
rect 25962 0 26018 800
rect 26514 0 26570 800
rect 26974 0 27030 800
rect 27526 0 27582 800
rect 28078 0 28134 800
rect 28538 0 28594 800
rect 29090 0 29146 800
rect 29550 0 29606 800
rect 30102 0 30158 800
rect 30654 0 30710 800
rect 31114 0 31170 800
rect 31666 0 31722 800
rect 32126 0 32182 800
rect 32678 0 32734 800
rect 33230 0 33286 800
rect 33690 0 33746 800
rect 34242 0 34298 800
rect 34794 0 34850 800
rect 35254 0 35310 800
rect 35806 0 35862 800
rect 36266 0 36322 800
rect 36818 0 36874 800
rect 37370 0 37426 800
rect 37830 0 37886 800
rect 38382 0 38438 800
rect 38842 0 38898 800
rect 39394 0 39450 800
rect 39946 0 40002 800
rect 40406 0 40462 800
rect 40958 0 41014 800
rect 41510 0 41566 800
rect 41970 0 42026 800
rect 42522 0 42578 800
rect 42982 0 43038 800
rect 43534 0 43590 800
rect 44086 0 44142 800
rect 44546 0 44602 800
rect 45098 0 45154 800
rect 45558 0 45614 800
rect 46110 0 46166 800
rect 46662 0 46718 800
rect 47122 0 47178 800
rect 47674 0 47730 800
rect 48134 0 48190 800
rect 48686 0 48742 800
rect 49238 0 49294 800
rect 49698 0 49754 800
rect 50250 0 50306 800
rect 50802 0 50858 800
rect 51262 0 51318 800
rect 51814 0 51870 800
rect 52274 0 52330 800
rect 52826 0 52882 800
rect 53378 0 53434 800
rect 53838 0 53894 800
rect 54390 0 54446 800
rect 54850 0 54906 800
rect 55402 0 55458 800
rect 55954 0 56010 800
rect 56414 0 56470 800
rect 56966 0 57022 800
rect 57426 0 57482 800
rect 57978 0 58034 800
rect 58530 0 58586 800
rect 58990 0 59046 800
rect 59542 0 59598 800
rect 60094 0 60150 800
rect 60554 0 60610 800
rect 61106 0 61162 800
rect 61566 0 61622 800
rect 62118 0 62174 800
rect 62670 0 62726 800
rect 63130 0 63186 800
rect 63682 0 63738 800
rect 64142 0 64198 800
rect 64694 0 64750 800
rect 65246 0 65302 800
rect 65706 0 65762 800
rect 66258 0 66314 800
rect 66810 0 66866 800
rect 67270 0 67326 800
rect 67822 0 67878 800
rect 68282 0 68338 800
rect 68834 0 68890 800
rect 69386 0 69442 800
rect 69846 0 69902 800
rect 70398 0 70454 800
rect 70858 0 70914 800
rect 71410 0 71466 800
rect 71962 0 72018 800
rect 72422 0 72478 800
rect 72974 0 73030 800
rect 73434 0 73490 800
rect 73986 0 74042 800
rect 74538 0 74594 800
rect 74998 0 75054 800
rect 75550 0 75606 800
rect 76102 0 76158 800
rect 76562 0 76618 800
rect 77114 0 77170 800
rect 77574 0 77630 800
rect 78126 0 78182 800
rect 78678 0 78734 800
rect 79138 0 79194 800
rect 79690 0 79746 800
rect 80150 0 80206 800
rect 80702 0 80758 800
rect 81254 0 81310 800
rect 81714 0 81770 800
rect 82266 0 82322 800
rect 82818 0 82874 800
rect 83278 0 83334 800
rect 83830 0 83886 800
rect 84290 0 84346 800
rect 84842 0 84898 800
rect 85394 0 85450 800
rect 85854 0 85910 800
rect 86406 0 86462 800
rect 86866 0 86922 800
rect 87418 0 87474 800
rect 87970 0 88026 800
rect 88430 0 88486 800
rect 88982 0 89038 800
rect 89442 0 89498 800
rect 89994 0 90050 800
rect 90546 0 90602 800
rect 91006 0 91062 800
rect 91558 0 91614 800
rect 92110 0 92166 800
rect 92570 0 92626 800
rect 93122 0 93178 800
rect 93582 0 93638 800
rect 94134 0 94190 800
rect 94686 0 94742 800
rect 95146 0 95202 800
rect 95698 0 95754 800
rect 96158 0 96214 800
rect 96710 0 96766 800
rect 97262 0 97318 800
rect 97722 0 97778 800
rect 98274 0 98330 800
rect 98826 0 98882 800
rect 99286 0 99342 800
rect 99838 0 99894 800
rect 100298 0 100354 800
rect 100850 0 100906 800
rect 101402 0 101458 800
rect 101862 0 101918 800
rect 102414 0 102470 800
rect 102874 0 102930 800
rect 103426 0 103482 800
rect 103978 0 104034 800
rect 104438 0 104494 800
rect 104990 0 105046 800
rect 105450 0 105506 800
rect 106002 0 106058 800
rect 106554 0 106610 800
rect 107014 0 107070 800
rect 107566 0 107622 800
rect 108118 0 108174 800
rect 108578 0 108634 800
rect 109130 0 109186 800
rect 109590 0 109646 800
rect 110142 0 110198 800
rect 110694 0 110750 800
rect 111154 0 111210 800
rect 111706 0 111762 800
rect 112166 0 112222 800
rect 112718 0 112774 800
rect 113270 0 113326 800
rect 113730 0 113786 800
rect 114282 0 114338 800
rect 114742 0 114798 800
rect 115294 0 115350 800
rect 115846 0 115902 800
rect 116306 0 116362 800
rect 116858 0 116914 800
rect 117410 0 117466 800
rect 117870 0 117926 800
rect 118422 0 118478 800
rect 118882 0 118938 800
rect 119434 0 119490 800
rect 119986 0 120042 800
rect 120446 0 120502 800
rect 120998 0 121054 800
rect 121458 0 121514 800
rect 122010 0 122066 800
rect 122562 0 122618 800
rect 123022 0 123078 800
rect 123574 0 123630 800
rect 124126 0 124182 800
rect 124586 0 124642 800
rect 125138 0 125194 800
rect 125598 0 125654 800
rect 126150 0 126206 800
rect 126702 0 126758 800
rect 127162 0 127218 800
rect 127714 0 127770 800
rect 128174 0 128230 800
rect 128726 0 128782 800
rect 129278 0 129334 800
rect 129738 0 129794 800
rect 130290 0 130346 800
rect 130750 0 130806 800
rect 131302 0 131358 800
rect 131854 0 131910 800
rect 132314 0 132370 800
rect 132866 0 132922 800
rect 133418 0 133474 800
rect 133878 0 133934 800
rect 134430 0 134486 800
rect 134890 0 134946 800
rect 135442 0 135498 800
rect 135994 0 136050 800
rect 136454 0 136510 800
rect 137006 0 137062 800
rect 137466 0 137522 800
rect 138018 0 138074 800
rect 138570 0 138626 800
rect 139030 0 139086 800
rect 139582 0 139638 800
rect 140134 0 140190 800
rect 140594 0 140650 800
rect 141146 0 141202 800
rect 141606 0 141662 800
rect 142158 0 142214 800
rect 142710 0 142766 800
rect 143170 0 143226 800
rect 143722 0 143778 800
rect 144182 0 144238 800
rect 144734 0 144790 800
rect 145286 0 145342 800
rect 145746 0 145802 800
rect 146298 0 146354 800
rect 146758 0 146814 800
rect 147310 0 147366 800
rect 147862 0 147918 800
rect 148322 0 148378 800
rect 148874 0 148930 800
rect 149426 0 149482 800
rect 149886 0 149942 800
rect 150438 0 150494 800
rect 150898 0 150954 800
rect 151450 0 151506 800
rect 152002 0 152058 800
rect 152462 0 152518 800
rect 153014 0 153070 800
rect 153474 0 153530 800
rect 154026 0 154082 800
rect 154578 0 154634 800
rect 155038 0 155094 800
rect 155590 0 155646 800
rect 156050 0 156106 800
rect 156602 0 156658 800
rect 157154 0 157210 800
rect 157614 0 157670 800
rect 158166 0 158222 800
rect 158718 0 158774 800
rect 159178 0 159234 800
rect 159730 0 159786 800
rect 160190 0 160246 800
rect 160742 0 160798 800
rect 161294 0 161350 800
rect 161754 0 161810 800
rect 162306 0 162362 800
rect 162766 0 162822 800
rect 163318 0 163374 800
rect 163870 0 163926 800
rect 164330 0 164386 800
rect 164882 0 164938 800
rect 165434 0 165490 800
rect 165894 0 165950 800
rect 166446 0 166502 800
rect 166906 0 166962 800
rect 167458 0 167514 800
rect 168010 0 168066 800
rect 168470 0 168526 800
rect 169022 0 169078 800
rect 169482 0 169538 800
rect 170034 0 170090 800
rect 170586 0 170642 800
rect 171046 0 171102 800
rect 171598 0 171654 800
rect 172058 0 172114 800
rect 172610 0 172666 800
rect 173162 0 173218 800
rect 173622 0 173678 800
rect 174174 0 174230 800
rect 174726 0 174782 800
rect 175186 0 175242 800
rect 175738 0 175794 800
rect 176198 0 176254 800
rect 176750 0 176806 800
rect 177302 0 177358 800
rect 177762 0 177818 800
rect 178314 0 178370 800
rect 178774 0 178830 800
rect 179326 0 179382 800
rect 179878 0 179934 800
rect 180338 0 180394 800
rect 180890 0 180946 800
rect 181442 0 181498 800
rect 181902 0 181958 800
rect 182454 0 182510 800
rect 182914 0 182970 800
rect 183466 0 183522 800
rect 184018 0 184074 800
rect 184478 0 184534 800
rect 185030 0 185086 800
rect 185490 0 185546 800
rect 186042 0 186098 800
rect 186594 0 186650 800
rect 187054 0 187110 800
rect 187606 0 187662 800
rect 188066 0 188122 800
rect 188618 0 188674 800
rect 189170 0 189226 800
rect 189630 0 189686 800
rect 190182 0 190238 800
rect 190734 0 190790 800
rect 191194 0 191250 800
rect 191746 0 191802 800
rect 192206 0 192262 800
rect 192758 0 192814 800
rect 193310 0 193366 800
rect 193770 0 193826 800
rect 194322 0 194378 800
rect 194782 0 194838 800
rect 195334 0 195390 800
rect 195886 0 195942 800
rect 196346 0 196402 800
rect 196898 0 196954 800
rect 197450 0 197506 800
rect 197910 0 197966 800
rect 198462 0 198518 800
rect 198922 0 198978 800
rect 199474 0 199530 800
rect 200026 0 200082 800
rect 200486 0 200542 800
rect 201038 0 201094 800
rect 201498 0 201554 800
rect 202050 0 202106 800
rect 202602 0 202658 800
rect 203062 0 203118 800
rect 203614 0 203670 800
rect 204074 0 204130 800
rect 204626 0 204682 800
rect 205178 0 205234 800
rect 205638 0 205694 800
rect 206190 0 206246 800
rect 206742 0 206798 800
rect 207202 0 207258 800
rect 207754 0 207810 800
rect 208214 0 208270 800
rect 208766 0 208822 800
rect 209318 0 209374 800
rect 209778 0 209834 800
rect 210330 0 210386 800
rect 210790 0 210846 800
rect 211342 0 211398 800
rect 211894 0 211950 800
rect 212354 0 212410 800
rect 212906 0 212962 800
rect 213366 0 213422 800
rect 213918 0 213974 800
rect 214470 0 214526 800
rect 214930 0 214986 800
rect 215482 0 215538 800
rect 216034 0 216090 800
rect 216494 0 216550 800
rect 217046 0 217102 800
rect 217506 0 217562 800
rect 218058 0 218114 800
rect 218610 0 218666 800
rect 219070 0 219126 800
rect 219622 0 219678 800
rect 220082 0 220138 800
rect 220634 0 220690 800
rect 221186 0 221242 800
rect 221646 0 221702 800
rect 222198 0 222254 800
rect 222750 0 222806 800
rect 223210 0 223266 800
rect 223762 0 223818 800
rect 224222 0 224278 800
rect 224774 0 224830 800
rect 225326 0 225382 800
rect 225786 0 225842 800
rect 226338 0 226394 800
rect 226798 0 226854 800
rect 227350 0 227406 800
rect 227902 0 227958 800
rect 228362 0 228418 800
rect 228914 0 228970 800
rect 229374 0 229430 800
rect 229926 0 229982 800
rect 230478 0 230534 800
rect 230938 0 230994 800
rect 231490 0 231546 800
rect 232042 0 232098 800
rect 232502 0 232558 800
rect 233054 0 233110 800
rect 233514 0 233570 800
rect 234066 0 234122 800
rect 234618 0 234674 800
rect 235078 0 235134 800
rect 235630 0 235686 800
rect 236090 0 236146 800
rect 236642 0 236698 800
rect 237194 0 237250 800
rect 237654 0 237710 800
rect 238206 0 238262 800
rect 238758 0 238814 800
rect 239218 0 239274 800
rect 239770 0 239826 800
rect 240230 0 240286 800
rect 240782 0 240838 800
rect 241334 0 241390 800
rect 241794 0 241850 800
rect 242346 0 242402 800
rect 242806 0 242862 800
rect 243358 0 243414 800
rect 243910 0 243966 800
rect 244370 0 244426 800
rect 244922 0 244978 800
rect 245382 0 245438 800
rect 245934 0 245990 800
rect 246486 0 246542 800
rect 246946 0 247002 800
rect 247498 0 247554 800
rect 248050 0 248106 800
rect 248510 0 248566 800
rect 249062 0 249118 800
rect 249522 0 249578 800
rect 250074 0 250130 800
rect 250626 0 250682 800
rect 251086 0 251142 800
rect 251638 0 251694 800
rect 252098 0 252154 800
rect 252650 0 252706 800
rect 253202 0 253258 800
rect 253662 0 253718 800
rect 254214 0 254270 800
<< obsm2 >>
rect 204 306283 1066 306354
rect 1234 306283 3274 306354
rect 3442 306283 5482 306354
rect 5650 306283 7690 306354
rect 7858 306283 9990 306354
rect 10158 306283 12198 306354
rect 12366 306283 14406 306354
rect 14574 306283 16614 306354
rect 16782 306283 18914 306354
rect 19082 306283 21122 306354
rect 21290 306283 23330 306354
rect 23498 306283 25538 306354
rect 25706 306283 27838 306354
rect 28006 306283 30046 306354
rect 30214 306283 32254 306354
rect 32422 306283 34554 306354
rect 34722 306283 36762 306354
rect 36930 306283 38970 306354
rect 39138 306283 41178 306354
rect 41346 306283 43478 306354
rect 43646 306283 45686 306354
rect 45854 306283 47894 306354
rect 48062 306283 50102 306354
rect 50270 306283 52402 306354
rect 52570 306283 54610 306354
rect 54778 306283 56818 306354
rect 56986 306283 59118 306354
rect 59286 306283 61326 306354
rect 61494 306283 63534 306354
rect 63702 306283 65742 306354
rect 65910 306283 68042 306354
rect 68210 306283 70250 306354
rect 70418 306283 72458 306354
rect 72626 306283 74666 306354
rect 74834 306283 76966 306354
rect 77134 306283 79174 306354
rect 79342 306283 81382 306354
rect 81550 306283 83682 306354
rect 83850 306283 85890 306354
rect 86058 306283 88098 306354
rect 88266 306283 90306 306354
rect 90474 306283 92606 306354
rect 92774 306283 94814 306354
rect 94982 306283 97022 306354
rect 97190 306283 99230 306354
rect 99398 306283 101530 306354
rect 101698 306283 103738 306354
rect 103906 306283 105946 306354
rect 106114 306283 108246 306354
rect 108414 306283 110454 306354
rect 110622 306283 112662 306354
rect 112830 306283 114870 306354
rect 115038 306283 117170 306354
rect 117338 306283 119378 306354
rect 119546 306283 121586 306354
rect 121754 306283 123794 306354
rect 123962 306283 126094 306354
rect 126262 306283 128302 306354
rect 128470 306283 130510 306354
rect 130678 306283 132810 306354
rect 132978 306283 135018 306354
rect 135186 306283 137226 306354
rect 137394 306283 139434 306354
rect 139602 306283 141734 306354
rect 141902 306283 143942 306354
rect 144110 306283 146150 306354
rect 146318 306283 148358 306354
rect 148526 306283 150658 306354
rect 150826 306283 152866 306354
rect 153034 306283 155074 306354
rect 155242 306283 157374 306354
rect 157542 306283 159582 306354
rect 159750 306283 161790 306354
rect 161958 306283 163998 306354
rect 164166 306283 166298 306354
rect 166466 306283 168506 306354
rect 168674 306283 170714 306354
rect 170882 306283 172922 306354
rect 173090 306283 175222 306354
rect 175390 306283 177430 306354
rect 177598 306283 179638 306354
rect 179806 306283 181938 306354
rect 182106 306283 184146 306354
rect 184314 306283 186354 306354
rect 186522 306283 188562 306354
rect 188730 306283 190862 306354
rect 191030 306283 193070 306354
rect 193238 306283 195278 306354
rect 195446 306283 197486 306354
rect 197654 306283 199786 306354
rect 199954 306283 201994 306354
rect 202162 306283 204202 306354
rect 204370 306283 206502 306354
rect 206670 306283 208710 306354
rect 208878 306283 210918 306354
rect 211086 306283 213126 306354
rect 213294 306283 215426 306354
rect 215594 306283 217634 306354
rect 217802 306283 219842 306354
rect 220010 306283 222050 306354
rect 222218 306283 224350 306354
rect 224518 306283 226558 306354
rect 226726 306283 228766 306354
rect 228934 306283 231066 306354
rect 231234 306283 233274 306354
rect 233442 306283 235482 306354
rect 235650 306283 237690 306354
rect 237858 306283 239990 306354
rect 240158 306283 242198 306354
rect 242366 306283 244406 306354
rect 244574 306283 246614 306354
rect 246782 306283 248914 306354
rect 249082 306283 251122 306354
rect 251290 306283 253330 306354
rect 253498 306283 254268 306354
rect 204 856 254268 306283
rect 314 734 606 856
rect 774 734 1158 856
rect 1326 734 1618 856
rect 1786 734 2170 856
rect 2338 734 2722 856
rect 2890 734 3182 856
rect 3350 734 3734 856
rect 3902 734 4194 856
rect 4362 734 4746 856
rect 4914 734 5298 856
rect 5466 734 5758 856
rect 5926 734 6310 856
rect 6478 734 6770 856
rect 6938 734 7322 856
rect 7490 734 7874 856
rect 8042 734 8334 856
rect 8502 734 8886 856
rect 9054 734 9438 856
rect 9606 734 9898 856
rect 10066 734 10450 856
rect 10618 734 10910 856
rect 11078 734 11462 856
rect 11630 734 12014 856
rect 12182 734 12474 856
rect 12642 734 13026 856
rect 13194 734 13486 856
rect 13654 734 14038 856
rect 14206 734 14590 856
rect 14758 734 15050 856
rect 15218 734 15602 856
rect 15770 734 16062 856
rect 16230 734 16614 856
rect 16782 734 17166 856
rect 17334 734 17626 856
rect 17794 734 18178 856
rect 18346 734 18730 856
rect 18898 734 19190 856
rect 19358 734 19742 856
rect 19910 734 20202 856
rect 20370 734 20754 856
rect 20922 734 21306 856
rect 21474 734 21766 856
rect 21934 734 22318 856
rect 22486 734 22778 856
rect 22946 734 23330 856
rect 23498 734 23882 856
rect 24050 734 24342 856
rect 24510 734 24894 856
rect 25062 734 25446 856
rect 25614 734 25906 856
rect 26074 734 26458 856
rect 26626 734 26918 856
rect 27086 734 27470 856
rect 27638 734 28022 856
rect 28190 734 28482 856
rect 28650 734 29034 856
rect 29202 734 29494 856
rect 29662 734 30046 856
rect 30214 734 30598 856
rect 30766 734 31058 856
rect 31226 734 31610 856
rect 31778 734 32070 856
rect 32238 734 32622 856
rect 32790 734 33174 856
rect 33342 734 33634 856
rect 33802 734 34186 856
rect 34354 734 34738 856
rect 34906 734 35198 856
rect 35366 734 35750 856
rect 35918 734 36210 856
rect 36378 734 36762 856
rect 36930 734 37314 856
rect 37482 734 37774 856
rect 37942 734 38326 856
rect 38494 734 38786 856
rect 38954 734 39338 856
rect 39506 734 39890 856
rect 40058 734 40350 856
rect 40518 734 40902 856
rect 41070 734 41454 856
rect 41622 734 41914 856
rect 42082 734 42466 856
rect 42634 734 42926 856
rect 43094 734 43478 856
rect 43646 734 44030 856
rect 44198 734 44490 856
rect 44658 734 45042 856
rect 45210 734 45502 856
rect 45670 734 46054 856
rect 46222 734 46606 856
rect 46774 734 47066 856
rect 47234 734 47618 856
rect 47786 734 48078 856
rect 48246 734 48630 856
rect 48798 734 49182 856
rect 49350 734 49642 856
rect 49810 734 50194 856
rect 50362 734 50746 856
rect 50914 734 51206 856
rect 51374 734 51758 856
rect 51926 734 52218 856
rect 52386 734 52770 856
rect 52938 734 53322 856
rect 53490 734 53782 856
rect 53950 734 54334 856
rect 54502 734 54794 856
rect 54962 734 55346 856
rect 55514 734 55898 856
rect 56066 734 56358 856
rect 56526 734 56910 856
rect 57078 734 57370 856
rect 57538 734 57922 856
rect 58090 734 58474 856
rect 58642 734 58934 856
rect 59102 734 59486 856
rect 59654 734 60038 856
rect 60206 734 60498 856
rect 60666 734 61050 856
rect 61218 734 61510 856
rect 61678 734 62062 856
rect 62230 734 62614 856
rect 62782 734 63074 856
rect 63242 734 63626 856
rect 63794 734 64086 856
rect 64254 734 64638 856
rect 64806 734 65190 856
rect 65358 734 65650 856
rect 65818 734 66202 856
rect 66370 734 66754 856
rect 66922 734 67214 856
rect 67382 734 67766 856
rect 67934 734 68226 856
rect 68394 734 68778 856
rect 68946 734 69330 856
rect 69498 734 69790 856
rect 69958 734 70342 856
rect 70510 734 70802 856
rect 70970 734 71354 856
rect 71522 734 71906 856
rect 72074 734 72366 856
rect 72534 734 72918 856
rect 73086 734 73378 856
rect 73546 734 73930 856
rect 74098 734 74482 856
rect 74650 734 74942 856
rect 75110 734 75494 856
rect 75662 734 76046 856
rect 76214 734 76506 856
rect 76674 734 77058 856
rect 77226 734 77518 856
rect 77686 734 78070 856
rect 78238 734 78622 856
rect 78790 734 79082 856
rect 79250 734 79634 856
rect 79802 734 80094 856
rect 80262 734 80646 856
rect 80814 734 81198 856
rect 81366 734 81658 856
rect 81826 734 82210 856
rect 82378 734 82762 856
rect 82930 734 83222 856
rect 83390 734 83774 856
rect 83942 734 84234 856
rect 84402 734 84786 856
rect 84954 734 85338 856
rect 85506 734 85798 856
rect 85966 734 86350 856
rect 86518 734 86810 856
rect 86978 734 87362 856
rect 87530 734 87914 856
rect 88082 734 88374 856
rect 88542 734 88926 856
rect 89094 734 89386 856
rect 89554 734 89938 856
rect 90106 734 90490 856
rect 90658 734 90950 856
rect 91118 734 91502 856
rect 91670 734 92054 856
rect 92222 734 92514 856
rect 92682 734 93066 856
rect 93234 734 93526 856
rect 93694 734 94078 856
rect 94246 734 94630 856
rect 94798 734 95090 856
rect 95258 734 95642 856
rect 95810 734 96102 856
rect 96270 734 96654 856
rect 96822 734 97206 856
rect 97374 734 97666 856
rect 97834 734 98218 856
rect 98386 734 98770 856
rect 98938 734 99230 856
rect 99398 734 99782 856
rect 99950 734 100242 856
rect 100410 734 100794 856
rect 100962 734 101346 856
rect 101514 734 101806 856
rect 101974 734 102358 856
rect 102526 734 102818 856
rect 102986 734 103370 856
rect 103538 734 103922 856
rect 104090 734 104382 856
rect 104550 734 104934 856
rect 105102 734 105394 856
rect 105562 734 105946 856
rect 106114 734 106498 856
rect 106666 734 106958 856
rect 107126 734 107510 856
rect 107678 734 108062 856
rect 108230 734 108522 856
rect 108690 734 109074 856
rect 109242 734 109534 856
rect 109702 734 110086 856
rect 110254 734 110638 856
rect 110806 734 111098 856
rect 111266 734 111650 856
rect 111818 734 112110 856
rect 112278 734 112662 856
rect 112830 734 113214 856
rect 113382 734 113674 856
rect 113842 734 114226 856
rect 114394 734 114686 856
rect 114854 734 115238 856
rect 115406 734 115790 856
rect 115958 734 116250 856
rect 116418 734 116802 856
rect 116970 734 117354 856
rect 117522 734 117814 856
rect 117982 734 118366 856
rect 118534 734 118826 856
rect 118994 734 119378 856
rect 119546 734 119930 856
rect 120098 734 120390 856
rect 120558 734 120942 856
rect 121110 734 121402 856
rect 121570 734 121954 856
rect 122122 734 122506 856
rect 122674 734 122966 856
rect 123134 734 123518 856
rect 123686 734 124070 856
rect 124238 734 124530 856
rect 124698 734 125082 856
rect 125250 734 125542 856
rect 125710 734 126094 856
rect 126262 734 126646 856
rect 126814 734 127106 856
rect 127274 734 127658 856
rect 127826 734 128118 856
rect 128286 734 128670 856
rect 128838 734 129222 856
rect 129390 734 129682 856
rect 129850 734 130234 856
rect 130402 734 130694 856
rect 130862 734 131246 856
rect 131414 734 131798 856
rect 131966 734 132258 856
rect 132426 734 132810 856
rect 132978 734 133362 856
rect 133530 734 133822 856
rect 133990 734 134374 856
rect 134542 734 134834 856
rect 135002 734 135386 856
rect 135554 734 135938 856
rect 136106 734 136398 856
rect 136566 734 136950 856
rect 137118 734 137410 856
rect 137578 734 137962 856
rect 138130 734 138514 856
rect 138682 734 138974 856
rect 139142 734 139526 856
rect 139694 734 140078 856
rect 140246 734 140538 856
rect 140706 734 141090 856
rect 141258 734 141550 856
rect 141718 734 142102 856
rect 142270 734 142654 856
rect 142822 734 143114 856
rect 143282 734 143666 856
rect 143834 734 144126 856
rect 144294 734 144678 856
rect 144846 734 145230 856
rect 145398 734 145690 856
rect 145858 734 146242 856
rect 146410 734 146702 856
rect 146870 734 147254 856
rect 147422 734 147806 856
rect 147974 734 148266 856
rect 148434 734 148818 856
rect 148986 734 149370 856
rect 149538 734 149830 856
rect 149998 734 150382 856
rect 150550 734 150842 856
rect 151010 734 151394 856
rect 151562 734 151946 856
rect 152114 734 152406 856
rect 152574 734 152958 856
rect 153126 734 153418 856
rect 153586 734 153970 856
rect 154138 734 154522 856
rect 154690 734 154982 856
rect 155150 734 155534 856
rect 155702 734 155994 856
rect 156162 734 156546 856
rect 156714 734 157098 856
rect 157266 734 157558 856
rect 157726 734 158110 856
rect 158278 734 158662 856
rect 158830 734 159122 856
rect 159290 734 159674 856
rect 159842 734 160134 856
rect 160302 734 160686 856
rect 160854 734 161238 856
rect 161406 734 161698 856
rect 161866 734 162250 856
rect 162418 734 162710 856
rect 162878 734 163262 856
rect 163430 734 163814 856
rect 163982 734 164274 856
rect 164442 734 164826 856
rect 164994 734 165378 856
rect 165546 734 165838 856
rect 166006 734 166390 856
rect 166558 734 166850 856
rect 167018 734 167402 856
rect 167570 734 167954 856
rect 168122 734 168414 856
rect 168582 734 168966 856
rect 169134 734 169426 856
rect 169594 734 169978 856
rect 170146 734 170530 856
rect 170698 734 170990 856
rect 171158 734 171542 856
rect 171710 734 172002 856
rect 172170 734 172554 856
rect 172722 734 173106 856
rect 173274 734 173566 856
rect 173734 734 174118 856
rect 174286 734 174670 856
rect 174838 734 175130 856
rect 175298 734 175682 856
rect 175850 734 176142 856
rect 176310 734 176694 856
rect 176862 734 177246 856
rect 177414 734 177706 856
rect 177874 734 178258 856
rect 178426 734 178718 856
rect 178886 734 179270 856
rect 179438 734 179822 856
rect 179990 734 180282 856
rect 180450 734 180834 856
rect 181002 734 181386 856
rect 181554 734 181846 856
rect 182014 734 182398 856
rect 182566 734 182858 856
rect 183026 734 183410 856
rect 183578 734 183962 856
rect 184130 734 184422 856
rect 184590 734 184974 856
rect 185142 734 185434 856
rect 185602 734 185986 856
rect 186154 734 186538 856
rect 186706 734 186998 856
rect 187166 734 187550 856
rect 187718 734 188010 856
rect 188178 734 188562 856
rect 188730 734 189114 856
rect 189282 734 189574 856
rect 189742 734 190126 856
rect 190294 734 190678 856
rect 190846 734 191138 856
rect 191306 734 191690 856
rect 191858 734 192150 856
rect 192318 734 192702 856
rect 192870 734 193254 856
rect 193422 734 193714 856
rect 193882 734 194266 856
rect 194434 734 194726 856
rect 194894 734 195278 856
rect 195446 734 195830 856
rect 195998 734 196290 856
rect 196458 734 196842 856
rect 197010 734 197394 856
rect 197562 734 197854 856
rect 198022 734 198406 856
rect 198574 734 198866 856
rect 199034 734 199418 856
rect 199586 734 199970 856
rect 200138 734 200430 856
rect 200598 734 200982 856
rect 201150 734 201442 856
rect 201610 734 201994 856
rect 202162 734 202546 856
rect 202714 734 203006 856
rect 203174 734 203558 856
rect 203726 734 204018 856
rect 204186 734 204570 856
rect 204738 734 205122 856
rect 205290 734 205582 856
rect 205750 734 206134 856
rect 206302 734 206686 856
rect 206854 734 207146 856
rect 207314 734 207698 856
rect 207866 734 208158 856
rect 208326 734 208710 856
rect 208878 734 209262 856
rect 209430 734 209722 856
rect 209890 734 210274 856
rect 210442 734 210734 856
rect 210902 734 211286 856
rect 211454 734 211838 856
rect 212006 734 212298 856
rect 212466 734 212850 856
rect 213018 734 213310 856
rect 213478 734 213862 856
rect 214030 734 214414 856
rect 214582 734 214874 856
rect 215042 734 215426 856
rect 215594 734 215978 856
rect 216146 734 216438 856
rect 216606 734 216990 856
rect 217158 734 217450 856
rect 217618 734 218002 856
rect 218170 734 218554 856
rect 218722 734 219014 856
rect 219182 734 219566 856
rect 219734 734 220026 856
rect 220194 734 220578 856
rect 220746 734 221130 856
rect 221298 734 221590 856
rect 221758 734 222142 856
rect 222310 734 222694 856
rect 222862 734 223154 856
rect 223322 734 223706 856
rect 223874 734 224166 856
rect 224334 734 224718 856
rect 224886 734 225270 856
rect 225438 734 225730 856
rect 225898 734 226282 856
rect 226450 734 226742 856
rect 226910 734 227294 856
rect 227462 734 227846 856
rect 228014 734 228306 856
rect 228474 734 228858 856
rect 229026 734 229318 856
rect 229486 734 229870 856
rect 230038 734 230422 856
rect 230590 734 230882 856
rect 231050 734 231434 856
rect 231602 734 231986 856
rect 232154 734 232446 856
rect 232614 734 232998 856
rect 233166 734 233458 856
rect 233626 734 234010 856
rect 234178 734 234562 856
rect 234730 734 235022 856
rect 235190 734 235574 856
rect 235742 734 236034 856
rect 236202 734 236586 856
rect 236754 734 237138 856
rect 237306 734 237598 856
rect 237766 734 238150 856
rect 238318 734 238702 856
rect 238870 734 239162 856
rect 239330 734 239714 856
rect 239882 734 240174 856
rect 240342 734 240726 856
rect 240894 734 241278 856
rect 241446 734 241738 856
rect 241906 734 242290 856
rect 242458 734 242750 856
rect 242918 734 243302 856
rect 243470 734 243854 856
rect 244022 734 244314 856
rect 244482 734 244866 856
rect 245034 734 245326 856
rect 245494 734 245878 856
rect 246046 734 246430 856
rect 246598 734 246890 856
rect 247058 734 247442 856
rect 247610 734 247994 856
rect 248162 734 248454 856
rect 248622 734 249006 856
rect 249174 734 249466 856
rect 249634 734 250018 856
rect 250186 734 250570 856
rect 250738 734 251030 856
rect 251198 734 251582 856
rect 251750 734 252042 856
rect 252210 734 252594 856
rect 252762 734 253146 856
rect 253314 734 253606 856
rect 253774 734 254158 856
<< obsm3 >>
rect 657 2143 252251 304673
<< metal4 >>
rect 4208 2128 4528 304688
rect 19568 2128 19888 304688
rect 34928 2128 35248 304688
rect 50288 2128 50608 304688
rect 65648 2128 65968 304688
rect 81008 2128 81328 304688
rect 96368 2128 96688 304688
rect 111728 2128 112048 304688
rect 127088 2128 127408 304688
rect 142448 2128 142768 304688
rect 157808 2128 158128 304688
rect 173168 2128 173488 304688
rect 188528 2128 188848 304688
rect 203888 2128 204208 304688
rect 219248 2128 219568 304688
rect 234608 2128 234928 304688
rect 249968 2128 250288 304688
<< obsm4 >>
rect 3187 3027 4128 302293
rect 4608 3027 19488 302293
rect 19968 3027 34848 302293
rect 35328 3027 50208 302293
rect 50688 3027 65568 302293
rect 66048 3027 80928 302293
rect 81408 3027 96288 302293
rect 96768 3027 111648 302293
rect 112128 3027 127008 302293
rect 127488 3027 142368 302293
rect 142848 3027 157728 302293
rect 158208 3027 173088 302293
rect 173568 3027 188448 302293
rect 188928 3027 203808 302293
rect 204288 3027 219168 302293
rect 219648 3027 234528 302293
rect 235008 3027 249888 302293
rect 250368 3027 251101 302293
<< labels >>
rlabel metal2 s 1122 306339 1178 307139 6 io_in[0]
port 1 nsew signal input
rlabel metal2 s 68098 306339 68154 307139 6 io_in[10]
port 2 nsew signal input
rlabel metal2 s 74722 306339 74778 307139 6 io_in[11]
port 3 nsew signal input
rlabel metal2 s 81438 306339 81494 307139 6 io_in[12]
port 4 nsew signal input
rlabel metal2 s 88154 306339 88210 307139 6 io_in[13]
port 5 nsew signal input
rlabel metal2 s 94870 306339 94926 307139 6 io_in[14]
port 6 nsew signal input
rlabel metal2 s 101586 306339 101642 307139 6 io_in[15]
port 7 nsew signal input
rlabel metal2 s 108302 306339 108358 307139 6 io_in[16]
port 8 nsew signal input
rlabel metal2 s 114926 306339 114982 307139 6 io_in[17]
port 9 nsew signal input
rlabel metal2 s 121642 306339 121698 307139 6 io_in[18]
port 10 nsew signal input
rlabel metal2 s 128358 306339 128414 307139 6 io_in[19]
port 11 nsew signal input
rlabel metal2 s 7746 306339 7802 307139 6 io_in[1]
port 12 nsew signal input
rlabel metal2 s 135074 306339 135130 307139 6 io_in[20]
port 13 nsew signal input
rlabel metal2 s 141790 306339 141846 307139 6 io_in[21]
port 14 nsew signal input
rlabel metal2 s 148414 306339 148470 307139 6 io_in[22]
port 15 nsew signal input
rlabel metal2 s 155130 306339 155186 307139 6 io_in[23]
port 16 nsew signal input
rlabel metal2 s 161846 306339 161902 307139 6 io_in[24]
port 17 nsew signal input
rlabel metal2 s 168562 306339 168618 307139 6 io_in[25]
port 18 nsew signal input
rlabel metal2 s 175278 306339 175334 307139 6 io_in[26]
port 19 nsew signal input
rlabel metal2 s 181994 306339 182050 307139 6 io_in[27]
port 20 nsew signal input
rlabel metal2 s 188618 306339 188674 307139 6 io_in[28]
port 21 nsew signal input
rlabel metal2 s 195334 306339 195390 307139 6 io_in[29]
port 22 nsew signal input
rlabel metal2 s 14462 306339 14518 307139 6 io_in[2]
port 23 nsew signal input
rlabel metal2 s 202050 306339 202106 307139 6 io_in[30]
port 24 nsew signal input
rlabel metal2 s 208766 306339 208822 307139 6 io_in[31]
port 25 nsew signal input
rlabel metal2 s 215482 306339 215538 307139 6 io_in[32]
port 26 nsew signal input
rlabel metal2 s 222106 306339 222162 307139 6 io_in[33]
port 27 nsew signal input
rlabel metal2 s 228822 306339 228878 307139 6 io_in[34]
port 28 nsew signal input
rlabel metal2 s 235538 306339 235594 307139 6 io_in[35]
port 29 nsew signal input
rlabel metal2 s 242254 306339 242310 307139 6 io_in[36]
port 30 nsew signal input
rlabel metal2 s 248970 306339 249026 307139 6 io_in[37]
port 31 nsew signal input
rlabel metal2 s 21178 306339 21234 307139 6 io_in[3]
port 32 nsew signal input
rlabel metal2 s 27894 306339 27950 307139 6 io_in[4]
port 33 nsew signal input
rlabel metal2 s 34610 306339 34666 307139 6 io_in[5]
port 34 nsew signal input
rlabel metal2 s 41234 306339 41290 307139 6 io_in[6]
port 35 nsew signal input
rlabel metal2 s 47950 306339 48006 307139 6 io_in[7]
port 36 nsew signal input
rlabel metal2 s 54666 306339 54722 307139 6 io_in[8]
port 37 nsew signal input
rlabel metal2 s 61382 306339 61438 307139 6 io_in[9]
port 38 nsew signal input
rlabel metal2 s 3330 306339 3386 307139 6 io_oeb[0]
port 39 nsew signal output
rlabel metal2 s 70306 306339 70362 307139 6 io_oeb[10]
port 40 nsew signal output
rlabel metal2 s 77022 306339 77078 307139 6 io_oeb[11]
port 41 nsew signal output
rlabel metal2 s 83738 306339 83794 307139 6 io_oeb[12]
port 42 nsew signal output
rlabel metal2 s 90362 306339 90418 307139 6 io_oeb[13]
port 43 nsew signal output
rlabel metal2 s 97078 306339 97134 307139 6 io_oeb[14]
port 44 nsew signal output
rlabel metal2 s 103794 306339 103850 307139 6 io_oeb[15]
port 45 nsew signal output
rlabel metal2 s 110510 306339 110566 307139 6 io_oeb[16]
port 46 nsew signal output
rlabel metal2 s 117226 306339 117282 307139 6 io_oeb[17]
port 47 nsew signal output
rlabel metal2 s 123850 306339 123906 307139 6 io_oeb[18]
port 48 nsew signal output
rlabel metal2 s 130566 306339 130622 307139 6 io_oeb[19]
port 49 nsew signal output
rlabel metal2 s 10046 306339 10102 307139 6 io_oeb[1]
port 50 nsew signal output
rlabel metal2 s 137282 306339 137338 307139 6 io_oeb[20]
port 51 nsew signal output
rlabel metal2 s 143998 306339 144054 307139 6 io_oeb[21]
port 52 nsew signal output
rlabel metal2 s 150714 306339 150770 307139 6 io_oeb[22]
port 53 nsew signal output
rlabel metal2 s 157430 306339 157486 307139 6 io_oeb[23]
port 54 nsew signal output
rlabel metal2 s 164054 306339 164110 307139 6 io_oeb[24]
port 55 nsew signal output
rlabel metal2 s 170770 306339 170826 307139 6 io_oeb[25]
port 56 nsew signal output
rlabel metal2 s 177486 306339 177542 307139 6 io_oeb[26]
port 57 nsew signal output
rlabel metal2 s 184202 306339 184258 307139 6 io_oeb[27]
port 58 nsew signal output
rlabel metal2 s 190918 306339 190974 307139 6 io_oeb[28]
port 59 nsew signal output
rlabel metal2 s 197542 306339 197598 307139 6 io_oeb[29]
port 60 nsew signal output
rlabel metal2 s 16670 306339 16726 307139 6 io_oeb[2]
port 61 nsew signal output
rlabel metal2 s 204258 306339 204314 307139 6 io_oeb[30]
port 62 nsew signal output
rlabel metal2 s 210974 306339 211030 307139 6 io_oeb[31]
port 63 nsew signal output
rlabel metal2 s 217690 306339 217746 307139 6 io_oeb[32]
port 64 nsew signal output
rlabel metal2 s 224406 306339 224462 307139 6 io_oeb[33]
port 65 nsew signal output
rlabel metal2 s 231122 306339 231178 307139 6 io_oeb[34]
port 66 nsew signal output
rlabel metal2 s 237746 306339 237802 307139 6 io_oeb[35]
port 67 nsew signal output
rlabel metal2 s 244462 306339 244518 307139 6 io_oeb[36]
port 68 nsew signal output
rlabel metal2 s 251178 306339 251234 307139 6 io_oeb[37]
port 69 nsew signal output
rlabel metal2 s 23386 306339 23442 307139 6 io_oeb[3]
port 70 nsew signal output
rlabel metal2 s 30102 306339 30158 307139 6 io_oeb[4]
port 71 nsew signal output
rlabel metal2 s 36818 306339 36874 307139 6 io_oeb[5]
port 72 nsew signal output
rlabel metal2 s 43534 306339 43590 307139 6 io_oeb[6]
port 73 nsew signal output
rlabel metal2 s 50158 306339 50214 307139 6 io_oeb[7]
port 74 nsew signal output
rlabel metal2 s 56874 306339 56930 307139 6 io_oeb[8]
port 75 nsew signal output
rlabel metal2 s 63590 306339 63646 307139 6 io_oeb[9]
port 76 nsew signal output
rlabel metal2 s 5538 306339 5594 307139 6 io_out[0]
port 77 nsew signal output
rlabel metal2 s 72514 306339 72570 307139 6 io_out[10]
port 78 nsew signal output
rlabel metal2 s 79230 306339 79286 307139 6 io_out[11]
port 79 nsew signal output
rlabel metal2 s 85946 306339 86002 307139 6 io_out[12]
port 80 nsew signal output
rlabel metal2 s 92662 306339 92718 307139 6 io_out[13]
port 81 nsew signal output
rlabel metal2 s 99286 306339 99342 307139 6 io_out[14]
port 82 nsew signal output
rlabel metal2 s 106002 306339 106058 307139 6 io_out[15]
port 83 nsew signal output
rlabel metal2 s 112718 306339 112774 307139 6 io_out[16]
port 84 nsew signal output
rlabel metal2 s 119434 306339 119490 307139 6 io_out[17]
port 85 nsew signal output
rlabel metal2 s 126150 306339 126206 307139 6 io_out[18]
port 86 nsew signal output
rlabel metal2 s 132866 306339 132922 307139 6 io_out[19]
port 87 nsew signal output
rlabel metal2 s 12254 306339 12310 307139 6 io_out[1]
port 88 nsew signal output
rlabel metal2 s 139490 306339 139546 307139 6 io_out[20]
port 89 nsew signal output
rlabel metal2 s 146206 306339 146262 307139 6 io_out[21]
port 90 nsew signal output
rlabel metal2 s 152922 306339 152978 307139 6 io_out[22]
port 91 nsew signal output
rlabel metal2 s 159638 306339 159694 307139 6 io_out[23]
port 92 nsew signal output
rlabel metal2 s 166354 306339 166410 307139 6 io_out[24]
port 93 nsew signal output
rlabel metal2 s 172978 306339 173034 307139 6 io_out[25]
port 94 nsew signal output
rlabel metal2 s 179694 306339 179750 307139 6 io_out[26]
port 95 nsew signal output
rlabel metal2 s 186410 306339 186466 307139 6 io_out[27]
port 96 nsew signal output
rlabel metal2 s 193126 306339 193182 307139 6 io_out[28]
port 97 nsew signal output
rlabel metal2 s 199842 306339 199898 307139 6 io_out[29]
port 98 nsew signal output
rlabel metal2 s 18970 306339 19026 307139 6 io_out[2]
port 99 nsew signal output
rlabel metal2 s 206558 306339 206614 307139 6 io_out[30]
port 100 nsew signal output
rlabel metal2 s 213182 306339 213238 307139 6 io_out[31]
port 101 nsew signal output
rlabel metal2 s 219898 306339 219954 307139 6 io_out[32]
port 102 nsew signal output
rlabel metal2 s 226614 306339 226670 307139 6 io_out[33]
port 103 nsew signal output
rlabel metal2 s 233330 306339 233386 307139 6 io_out[34]
port 104 nsew signal output
rlabel metal2 s 240046 306339 240102 307139 6 io_out[35]
port 105 nsew signal output
rlabel metal2 s 246670 306339 246726 307139 6 io_out[36]
port 106 nsew signal output
rlabel metal2 s 253386 306339 253442 307139 6 io_out[37]
port 107 nsew signal output
rlabel metal2 s 25594 306339 25650 307139 6 io_out[3]
port 108 nsew signal output
rlabel metal2 s 32310 306339 32366 307139 6 io_out[4]
port 109 nsew signal output
rlabel metal2 s 39026 306339 39082 307139 6 io_out[5]
port 110 nsew signal output
rlabel metal2 s 45742 306339 45798 307139 6 io_out[6]
port 111 nsew signal output
rlabel metal2 s 52458 306339 52514 307139 6 io_out[7]
port 112 nsew signal output
rlabel metal2 s 59174 306339 59230 307139 6 io_out[8]
port 113 nsew signal output
rlabel metal2 s 65798 306339 65854 307139 6 io_out[9]
port 114 nsew signal output
rlabel metal2 s 253202 0 253258 800 6 irq[0]
port 115 nsew signal output
rlabel metal2 s 253662 0 253718 800 6 irq[1]
port 116 nsew signal output
rlabel metal2 s 254214 0 254270 800 6 irq[2]
port 117 nsew signal output
rlabel metal2 s 54850 0 54906 800 6 la_data_in[0]
port 118 nsew signal input
rlabel metal2 s 209778 0 209834 800 6 la_data_in[100]
port 119 nsew signal input
rlabel metal2 s 211342 0 211398 800 6 la_data_in[101]
port 120 nsew signal input
rlabel metal2 s 212906 0 212962 800 6 la_data_in[102]
port 121 nsew signal input
rlabel metal2 s 214470 0 214526 800 6 la_data_in[103]
port 122 nsew signal input
rlabel metal2 s 216034 0 216090 800 6 la_data_in[104]
port 123 nsew signal input
rlabel metal2 s 217506 0 217562 800 6 la_data_in[105]
port 124 nsew signal input
rlabel metal2 s 219070 0 219126 800 6 la_data_in[106]
port 125 nsew signal input
rlabel metal2 s 220634 0 220690 800 6 la_data_in[107]
port 126 nsew signal input
rlabel metal2 s 222198 0 222254 800 6 la_data_in[108]
port 127 nsew signal input
rlabel metal2 s 223762 0 223818 800 6 la_data_in[109]
port 128 nsew signal input
rlabel metal2 s 70398 0 70454 800 6 la_data_in[10]
port 129 nsew signal input
rlabel metal2 s 225326 0 225382 800 6 la_data_in[110]
port 130 nsew signal input
rlabel metal2 s 226798 0 226854 800 6 la_data_in[111]
port 131 nsew signal input
rlabel metal2 s 228362 0 228418 800 6 la_data_in[112]
port 132 nsew signal input
rlabel metal2 s 229926 0 229982 800 6 la_data_in[113]
port 133 nsew signal input
rlabel metal2 s 231490 0 231546 800 6 la_data_in[114]
port 134 nsew signal input
rlabel metal2 s 233054 0 233110 800 6 la_data_in[115]
port 135 nsew signal input
rlabel metal2 s 234618 0 234674 800 6 la_data_in[116]
port 136 nsew signal input
rlabel metal2 s 236090 0 236146 800 6 la_data_in[117]
port 137 nsew signal input
rlabel metal2 s 237654 0 237710 800 6 la_data_in[118]
port 138 nsew signal input
rlabel metal2 s 239218 0 239274 800 6 la_data_in[119]
port 139 nsew signal input
rlabel metal2 s 71962 0 72018 800 6 la_data_in[11]
port 140 nsew signal input
rlabel metal2 s 240782 0 240838 800 6 la_data_in[120]
port 141 nsew signal input
rlabel metal2 s 242346 0 242402 800 6 la_data_in[121]
port 142 nsew signal input
rlabel metal2 s 243910 0 243966 800 6 la_data_in[122]
port 143 nsew signal input
rlabel metal2 s 245382 0 245438 800 6 la_data_in[123]
port 144 nsew signal input
rlabel metal2 s 246946 0 247002 800 6 la_data_in[124]
port 145 nsew signal input
rlabel metal2 s 248510 0 248566 800 6 la_data_in[125]
port 146 nsew signal input
rlabel metal2 s 250074 0 250130 800 6 la_data_in[126]
port 147 nsew signal input
rlabel metal2 s 251638 0 251694 800 6 la_data_in[127]
port 148 nsew signal input
rlabel metal2 s 73434 0 73490 800 6 la_data_in[12]
port 149 nsew signal input
rlabel metal2 s 74998 0 75054 800 6 la_data_in[13]
port 150 nsew signal input
rlabel metal2 s 76562 0 76618 800 6 la_data_in[14]
port 151 nsew signal input
rlabel metal2 s 78126 0 78182 800 6 la_data_in[15]
port 152 nsew signal input
rlabel metal2 s 79690 0 79746 800 6 la_data_in[16]
port 153 nsew signal input
rlabel metal2 s 81254 0 81310 800 6 la_data_in[17]
port 154 nsew signal input
rlabel metal2 s 82818 0 82874 800 6 la_data_in[18]
port 155 nsew signal input
rlabel metal2 s 84290 0 84346 800 6 la_data_in[19]
port 156 nsew signal input
rlabel metal2 s 56414 0 56470 800 6 la_data_in[1]
port 157 nsew signal input
rlabel metal2 s 85854 0 85910 800 6 la_data_in[20]
port 158 nsew signal input
rlabel metal2 s 87418 0 87474 800 6 la_data_in[21]
port 159 nsew signal input
rlabel metal2 s 88982 0 89038 800 6 la_data_in[22]
port 160 nsew signal input
rlabel metal2 s 90546 0 90602 800 6 la_data_in[23]
port 161 nsew signal input
rlabel metal2 s 92110 0 92166 800 6 la_data_in[24]
port 162 nsew signal input
rlabel metal2 s 93582 0 93638 800 6 la_data_in[25]
port 163 nsew signal input
rlabel metal2 s 95146 0 95202 800 6 la_data_in[26]
port 164 nsew signal input
rlabel metal2 s 96710 0 96766 800 6 la_data_in[27]
port 165 nsew signal input
rlabel metal2 s 98274 0 98330 800 6 la_data_in[28]
port 166 nsew signal input
rlabel metal2 s 99838 0 99894 800 6 la_data_in[29]
port 167 nsew signal input
rlabel metal2 s 57978 0 58034 800 6 la_data_in[2]
port 168 nsew signal input
rlabel metal2 s 101402 0 101458 800 6 la_data_in[30]
port 169 nsew signal input
rlabel metal2 s 102874 0 102930 800 6 la_data_in[31]
port 170 nsew signal input
rlabel metal2 s 104438 0 104494 800 6 la_data_in[32]
port 171 nsew signal input
rlabel metal2 s 106002 0 106058 800 6 la_data_in[33]
port 172 nsew signal input
rlabel metal2 s 107566 0 107622 800 6 la_data_in[34]
port 173 nsew signal input
rlabel metal2 s 109130 0 109186 800 6 la_data_in[35]
port 174 nsew signal input
rlabel metal2 s 110694 0 110750 800 6 la_data_in[36]
port 175 nsew signal input
rlabel metal2 s 112166 0 112222 800 6 la_data_in[37]
port 176 nsew signal input
rlabel metal2 s 113730 0 113786 800 6 la_data_in[38]
port 177 nsew signal input
rlabel metal2 s 115294 0 115350 800 6 la_data_in[39]
port 178 nsew signal input
rlabel metal2 s 59542 0 59598 800 6 la_data_in[3]
port 179 nsew signal input
rlabel metal2 s 116858 0 116914 800 6 la_data_in[40]
port 180 nsew signal input
rlabel metal2 s 118422 0 118478 800 6 la_data_in[41]
port 181 nsew signal input
rlabel metal2 s 119986 0 120042 800 6 la_data_in[42]
port 182 nsew signal input
rlabel metal2 s 121458 0 121514 800 6 la_data_in[43]
port 183 nsew signal input
rlabel metal2 s 123022 0 123078 800 6 la_data_in[44]
port 184 nsew signal input
rlabel metal2 s 124586 0 124642 800 6 la_data_in[45]
port 185 nsew signal input
rlabel metal2 s 126150 0 126206 800 6 la_data_in[46]
port 186 nsew signal input
rlabel metal2 s 127714 0 127770 800 6 la_data_in[47]
port 187 nsew signal input
rlabel metal2 s 129278 0 129334 800 6 la_data_in[48]
port 188 nsew signal input
rlabel metal2 s 130750 0 130806 800 6 la_data_in[49]
port 189 nsew signal input
rlabel metal2 s 61106 0 61162 800 6 la_data_in[4]
port 190 nsew signal input
rlabel metal2 s 132314 0 132370 800 6 la_data_in[50]
port 191 nsew signal input
rlabel metal2 s 133878 0 133934 800 6 la_data_in[51]
port 192 nsew signal input
rlabel metal2 s 135442 0 135498 800 6 la_data_in[52]
port 193 nsew signal input
rlabel metal2 s 137006 0 137062 800 6 la_data_in[53]
port 194 nsew signal input
rlabel metal2 s 138570 0 138626 800 6 la_data_in[54]
port 195 nsew signal input
rlabel metal2 s 140134 0 140190 800 6 la_data_in[55]
port 196 nsew signal input
rlabel metal2 s 141606 0 141662 800 6 la_data_in[56]
port 197 nsew signal input
rlabel metal2 s 143170 0 143226 800 6 la_data_in[57]
port 198 nsew signal input
rlabel metal2 s 144734 0 144790 800 6 la_data_in[58]
port 199 nsew signal input
rlabel metal2 s 146298 0 146354 800 6 la_data_in[59]
port 200 nsew signal input
rlabel metal2 s 62670 0 62726 800 6 la_data_in[5]
port 201 nsew signal input
rlabel metal2 s 147862 0 147918 800 6 la_data_in[60]
port 202 nsew signal input
rlabel metal2 s 149426 0 149482 800 6 la_data_in[61]
port 203 nsew signal input
rlabel metal2 s 150898 0 150954 800 6 la_data_in[62]
port 204 nsew signal input
rlabel metal2 s 152462 0 152518 800 6 la_data_in[63]
port 205 nsew signal input
rlabel metal2 s 154026 0 154082 800 6 la_data_in[64]
port 206 nsew signal input
rlabel metal2 s 155590 0 155646 800 6 la_data_in[65]
port 207 nsew signal input
rlabel metal2 s 157154 0 157210 800 6 la_data_in[66]
port 208 nsew signal input
rlabel metal2 s 158718 0 158774 800 6 la_data_in[67]
port 209 nsew signal input
rlabel metal2 s 160190 0 160246 800 6 la_data_in[68]
port 210 nsew signal input
rlabel metal2 s 161754 0 161810 800 6 la_data_in[69]
port 211 nsew signal input
rlabel metal2 s 64142 0 64198 800 6 la_data_in[6]
port 212 nsew signal input
rlabel metal2 s 163318 0 163374 800 6 la_data_in[70]
port 213 nsew signal input
rlabel metal2 s 164882 0 164938 800 6 la_data_in[71]
port 214 nsew signal input
rlabel metal2 s 166446 0 166502 800 6 la_data_in[72]
port 215 nsew signal input
rlabel metal2 s 168010 0 168066 800 6 la_data_in[73]
port 216 nsew signal input
rlabel metal2 s 169482 0 169538 800 6 la_data_in[74]
port 217 nsew signal input
rlabel metal2 s 171046 0 171102 800 6 la_data_in[75]
port 218 nsew signal input
rlabel metal2 s 172610 0 172666 800 6 la_data_in[76]
port 219 nsew signal input
rlabel metal2 s 174174 0 174230 800 6 la_data_in[77]
port 220 nsew signal input
rlabel metal2 s 175738 0 175794 800 6 la_data_in[78]
port 221 nsew signal input
rlabel metal2 s 177302 0 177358 800 6 la_data_in[79]
port 222 nsew signal input
rlabel metal2 s 65706 0 65762 800 6 la_data_in[7]
port 223 nsew signal input
rlabel metal2 s 178774 0 178830 800 6 la_data_in[80]
port 224 nsew signal input
rlabel metal2 s 180338 0 180394 800 6 la_data_in[81]
port 225 nsew signal input
rlabel metal2 s 181902 0 181958 800 6 la_data_in[82]
port 226 nsew signal input
rlabel metal2 s 183466 0 183522 800 6 la_data_in[83]
port 227 nsew signal input
rlabel metal2 s 185030 0 185086 800 6 la_data_in[84]
port 228 nsew signal input
rlabel metal2 s 186594 0 186650 800 6 la_data_in[85]
port 229 nsew signal input
rlabel metal2 s 188066 0 188122 800 6 la_data_in[86]
port 230 nsew signal input
rlabel metal2 s 189630 0 189686 800 6 la_data_in[87]
port 231 nsew signal input
rlabel metal2 s 191194 0 191250 800 6 la_data_in[88]
port 232 nsew signal input
rlabel metal2 s 192758 0 192814 800 6 la_data_in[89]
port 233 nsew signal input
rlabel metal2 s 67270 0 67326 800 6 la_data_in[8]
port 234 nsew signal input
rlabel metal2 s 194322 0 194378 800 6 la_data_in[90]
port 235 nsew signal input
rlabel metal2 s 195886 0 195942 800 6 la_data_in[91]
port 236 nsew signal input
rlabel metal2 s 197450 0 197506 800 6 la_data_in[92]
port 237 nsew signal input
rlabel metal2 s 198922 0 198978 800 6 la_data_in[93]
port 238 nsew signal input
rlabel metal2 s 200486 0 200542 800 6 la_data_in[94]
port 239 nsew signal input
rlabel metal2 s 202050 0 202106 800 6 la_data_in[95]
port 240 nsew signal input
rlabel metal2 s 203614 0 203670 800 6 la_data_in[96]
port 241 nsew signal input
rlabel metal2 s 205178 0 205234 800 6 la_data_in[97]
port 242 nsew signal input
rlabel metal2 s 206742 0 206798 800 6 la_data_in[98]
port 243 nsew signal input
rlabel metal2 s 208214 0 208270 800 6 la_data_in[99]
port 244 nsew signal input
rlabel metal2 s 68834 0 68890 800 6 la_data_in[9]
port 245 nsew signal input
rlabel metal2 s 55402 0 55458 800 6 la_data_out[0]
port 246 nsew signal output
rlabel metal2 s 210330 0 210386 800 6 la_data_out[100]
port 247 nsew signal output
rlabel metal2 s 211894 0 211950 800 6 la_data_out[101]
port 248 nsew signal output
rlabel metal2 s 213366 0 213422 800 6 la_data_out[102]
port 249 nsew signal output
rlabel metal2 s 214930 0 214986 800 6 la_data_out[103]
port 250 nsew signal output
rlabel metal2 s 216494 0 216550 800 6 la_data_out[104]
port 251 nsew signal output
rlabel metal2 s 218058 0 218114 800 6 la_data_out[105]
port 252 nsew signal output
rlabel metal2 s 219622 0 219678 800 6 la_data_out[106]
port 253 nsew signal output
rlabel metal2 s 221186 0 221242 800 6 la_data_out[107]
port 254 nsew signal output
rlabel metal2 s 222750 0 222806 800 6 la_data_out[108]
port 255 nsew signal output
rlabel metal2 s 224222 0 224278 800 6 la_data_out[109]
port 256 nsew signal output
rlabel metal2 s 70858 0 70914 800 6 la_data_out[10]
port 257 nsew signal output
rlabel metal2 s 225786 0 225842 800 6 la_data_out[110]
port 258 nsew signal output
rlabel metal2 s 227350 0 227406 800 6 la_data_out[111]
port 259 nsew signal output
rlabel metal2 s 228914 0 228970 800 6 la_data_out[112]
port 260 nsew signal output
rlabel metal2 s 230478 0 230534 800 6 la_data_out[113]
port 261 nsew signal output
rlabel metal2 s 232042 0 232098 800 6 la_data_out[114]
port 262 nsew signal output
rlabel metal2 s 233514 0 233570 800 6 la_data_out[115]
port 263 nsew signal output
rlabel metal2 s 235078 0 235134 800 6 la_data_out[116]
port 264 nsew signal output
rlabel metal2 s 236642 0 236698 800 6 la_data_out[117]
port 265 nsew signal output
rlabel metal2 s 238206 0 238262 800 6 la_data_out[118]
port 266 nsew signal output
rlabel metal2 s 239770 0 239826 800 6 la_data_out[119]
port 267 nsew signal output
rlabel metal2 s 72422 0 72478 800 6 la_data_out[11]
port 268 nsew signal output
rlabel metal2 s 241334 0 241390 800 6 la_data_out[120]
port 269 nsew signal output
rlabel metal2 s 242806 0 242862 800 6 la_data_out[121]
port 270 nsew signal output
rlabel metal2 s 244370 0 244426 800 6 la_data_out[122]
port 271 nsew signal output
rlabel metal2 s 245934 0 245990 800 6 la_data_out[123]
port 272 nsew signal output
rlabel metal2 s 247498 0 247554 800 6 la_data_out[124]
port 273 nsew signal output
rlabel metal2 s 249062 0 249118 800 6 la_data_out[125]
port 274 nsew signal output
rlabel metal2 s 250626 0 250682 800 6 la_data_out[126]
port 275 nsew signal output
rlabel metal2 s 252098 0 252154 800 6 la_data_out[127]
port 276 nsew signal output
rlabel metal2 s 73986 0 74042 800 6 la_data_out[12]
port 277 nsew signal output
rlabel metal2 s 75550 0 75606 800 6 la_data_out[13]
port 278 nsew signal output
rlabel metal2 s 77114 0 77170 800 6 la_data_out[14]
port 279 nsew signal output
rlabel metal2 s 78678 0 78734 800 6 la_data_out[15]
port 280 nsew signal output
rlabel metal2 s 80150 0 80206 800 6 la_data_out[16]
port 281 nsew signal output
rlabel metal2 s 81714 0 81770 800 6 la_data_out[17]
port 282 nsew signal output
rlabel metal2 s 83278 0 83334 800 6 la_data_out[18]
port 283 nsew signal output
rlabel metal2 s 84842 0 84898 800 6 la_data_out[19]
port 284 nsew signal output
rlabel metal2 s 56966 0 57022 800 6 la_data_out[1]
port 285 nsew signal output
rlabel metal2 s 86406 0 86462 800 6 la_data_out[20]
port 286 nsew signal output
rlabel metal2 s 87970 0 88026 800 6 la_data_out[21]
port 287 nsew signal output
rlabel metal2 s 89442 0 89498 800 6 la_data_out[22]
port 288 nsew signal output
rlabel metal2 s 91006 0 91062 800 6 la_data_out[23]
port 289 nsew signal output
rlabel metal2 s 92570 0 92626 800 6 la_data_out[24]
port 290 nsew signal output
rlabel metal2 s 94134 0 94190 800 6 la_data_out[25]
port 291 nsew signal output
rlabel metal2 s 95698 0 95754 800 6 la_data_out[26]
port 292 nsew signal output
rlabel metal2 s 97262 0 97318 800 6 la_data_out[27]
port 293 nsew signal output
rlabel metal2 s 98826 0 98882 800 6 la_data_out[28]
port 294 nsew signal output
rlabel metal2 s 100298 0 100354 800 6 la_data_out[29]
port 295 nsew signal output
rlabel metal2 s 58530 0 58586 800 6 la_data_out[2]
port 296 nsew signal output
rlabel metal2 s 101862 0 101918 800 6 la_data_out[30]
port 297 nsew signal output
rlabel metal2 s 103426 0 103482 800 6 la_data_out[31]
port 298 nsew signal output
rlabel metal2 s 104990 0 105046 800 6 la_data_out[32]
port 299 nsew signal output
rlabel metal2 s 106554 0 106610 800 6 la_data_out[33]
port 300 nsew signal output
rlabel metal2 s 108118 0 108174 800 6 la_data_out[34]
port 301 nsew signal output
rlabel metal2 s 109590 0 109646 800 6 la_data_out[35]
port 302 nsew signal output
rlabel metal2 s 111154 0 111210 800 6 la_data_out[36]
port 303 nsew signal output
rlabel metal2 s 112718 0 112774 800 6 la_data_out[37]
port 304 nsew signal output
rlabel metal2 s 114282 0 114338 800 6 la_data_out[38]
port 305 nsew signal output
rlabel metal2 s 115846 0 115902 800 6 la_data_out[39]
port 306 nsew signal output
rlabel metal2 s 60094 0 60150 800 6 la_data_out[3]
port 307 nsew signal output
rlabel metal2 s 117410 0 117466 800 6 la_data_out[40]
port 308 nsew signal output
rlabel metal2 s 118882 0 118938 800 6 la_data_out[41]
port 309 nsew signal output
rlabel metal2 s 120446 0 120502 800 6 la_data_out[42]
port 310 nsew signal output
rlabel metal2 s 122010 0 122066 800 6 la_data_out[43]
port 311 nsew signal output
rlabel metal2 s 123574 0 123630 800 6 la_data_out[44]
port 312 nsew signal output
rlabel metal2 s 125138 0 125194 800 6 la_data_out[45]
port 313 nsew signal output
rlabel metal2 s 126702 0 126758 800 6 la_data_out[46]
port 314 nsew signal output
rlabel metal2 s 128174 0 128230 800 6 la_data_out[47]
port 315 nsew signal output
rlabel metal2 s 129738 0 129794 800 6 la_data_out[48]
port 316 nsew signal output
rlabel metal2 s 131302 0 131358 800 6 la_data_out[49]
port 317 nsew signal output
rlabel metal2 s 61566 0 61622 800 6 la_data_out[4]
port 318 nsew signal output
rlabel metal2 s 132866 0 132922 800 6 la_data_out[50]
port 319 nsew signal output
rlabel metal2 s 134430 0 134486 800 6 la_data_out[51]
port 320 nsew signal output
rlabel metal2 s 135994 0 136050 800 6 la_data_out[52]
port 321 nsew signal output
rlabel metal2 s 137466 0 137522 800 6 la_data_out[53]
port 322 nsew signal output
rlabel metal2 s 139030 0 139086 800 6 la_data_out[54]
port 323 nsew signal output
rlabel metal2 s 140594 0 140650 800 6 la_data_out[55]
port 324 nsew signal output
rlabel metal2 s 142158 0 142214 800 6 la_data_out[56]
port 325 nsew signal output
rlabel metal2 s 143722 0 143778 800 6 la_data_out[57]
port 326 nsew signal output
rlabel metal2 s 145286 0 145342 800 6 la_data_out[58]
port 327 nsew signal output
rlabel metal2 s 146758 0 146814 800 6 la_data_out[59]
port 328 nsew signal output
rlabel metal2 s 63130 0 63186 800 6 la_data_out[5]
port 329 nsew signal output
rlabel metal2 s 148322 0 148378 800 6 la_data_out[60]
port 330 nsew signal output
rlabel metal2 s 149886 0 149942 800 6 la_data_out[61]
port 331 nsew signal output
rlabel metal2 s 151450 0 151506 800 6 la_data_out[62]
port 332 nsew signal output
rlabel metal2 s 153014 0 153070 800 6 la_data_out[63]
port 333 nsew signal output
rlabel metal2 s 154578 0 154634 800 6 la_data_out[64]
port 334 nsew signal output
rlabel metal2 s 156050 0 156106 800 6 la_data_out[65]
port 335 nsew signal output
rlabel metal2 s 157614 0 157670 800 6 la_data_out[66]
port 336 nsew signal output
rlabel metal2 s 159178 0 159234 800 6 la_data_out[67]
port 337 nsew signal output
rlabel metal2 s 160742 0 160798 800 6 la_data_out[68]
port 338 nsew signal output
rlabel metal2 s 162306 0 162362 800 6 la_data_out[69]
port 339 nsew signal output
rlabel metal2 s 64694 0 64750 800 6 la_data_out[6]
port 340 nsew signal output
rlabel metal2 s 163870 0 163926 800 6 la_data_out[70]
port 341 nsew signal output
rlabel metal2 s 165434 0 165490 800 6 la_data_out[71]
port 342 nsew signal output
rlabel metal2 s 166906 0 166962 800 6 la_data_out[72]
port 343 nsew signal output
rlabel metal2 s 168470 0 168526 800 6 la_data_out[73]
port 344 nsew signal output
rlabel metal2 s 170034 0 170090 800 6 la_data_out[74]
port 345 nsew signal output
rlabel metal2 s 171598 0 171654 800 6 la_data_out[75]
port 346 nsew signal output
rlabel metal2 s 173162 0 173218 800 6 la_data_out[76]
port 347 nsew signal output
rlabel metal2 s 174726 0 174782 800 6 la_data_out[77]
port 348 nsew signal output
rlabel metal2 s 176198 0 176254 800 6 la_data_out[78]
port 349 nsew signal output
rlabel metal2 s 177762 0 177818 800 6 la_data_out[79]
port 350 nsew signal output
rlabel metal2 s 66258 0 66314 800 6 la_data_out[7]
port 351 nsew signal output
rlabel metal2 s 179326 0 179382 800 6 la_data_out[80]
port 352 nsew signal output
rlabel metal2 s 180890 0 180946 800 6 la_data_out[81]
port 353 nsew signal output
rlabel metal2 s 182454 0 182510 800 6 la_data_out[82]
port 354 nsew signal output
rlabel metal2 s 184018 0 184074 800 6 la_data_out[83]
port 355 nsew signal output
rlabel metal2 s 185490 0 185546 800 6 la_data_out[84]
port 356 nsew signal output
rlabel metal2 s 187054 0 187110 800 6 la_data_out[85]
port 357 nsew signal output
rlabel metal2 s 188618 0 188674 800 6 la_data_out[86]
port 358 nsew signal output
rlabel metal2 s 190182 0 190238 800 6 la_data_out[87]
port 359 nsew signal output
rlabel metal2 s 191746 0 191802 800 6 la_data_out[88]
port 360 nsew signal output
rlabel metal2 s 193310 0 193366 800 6 la_data_out[89]
port 361 nsew signal output
rlabel metal2 s 67822 0 67878 800 6 la_data_out[8]
port 362 nsew signal output
rlabel metal2 s 194782 0 194838 800 6 la_data_out[90]
port 363 nsew signal output
rlabel metal2 s 196346 0 196402 800 6 la_data_out[91]
port 364 nsew signal output
rlabel metal2 s 197910 0 197966 800 6 la_data_out[92]
port 365 nsew signal output
rlabel metal2 s 199474 0 199530 800 6 la_data_out[93]
port 366 nsew signal output
rlabel metal2 s 201038 0 201094 800 6 la_data_out[94]
port 367 nsew signal output
rlabel metal2 s 202602 0 202658 800 6 la_data_out[95]
port 368 nsew signal output
rlabel metal2 s 204074 0 204130 800 6 la_data_out[96]
port 369 nsew signal output
rlabel metal2 s 205638 0 205694 800 6 la_data_out[97]
port 370 nsew signal output
rlabel metal2 s 207202 0 207258 800 6 la_data_out[98]
port 371 nsew signal output
rlabel metal2 s 208766 0 208822 800 6 la_data_out[99]
port 372 nsew signal output
rlabel metal2 s 69386 0 69442 800 6 la_data_out[9]
port 373 nsew signal output
rlabel metal2 s 55954 0 56010 800 6 la_oenb[0]
port 374 nsew signal input
rlabel metal2 s 210790 0 210846 800 6 la_oenb[100]
port 375 nsew signal input
rlabel metal2 s 212354 0 212410 800 6 la_oenb[101]
port 376 nsew signal input
rlabel metal2 s 213918 0 213974 800 6 la_oenb[102]
port 377 nsew signal input
rlabel metal2 s 215482 0 215538 800 6 la_oenb[103]
port 378 nsew signal input
rlabel metal2 s 217046 0 217102 800 6 la_oenb[104]
port 379 nsew signal input
rlabel metal2 s 218610 0 218666 800 6 la_oenb[105]
port 380 nsew signal input
rlabel metal2 s 220082 0 220138 800 6 la_oenb[106]
port 381 nsew signal input
rlabel metal2 s 221646 0 221702 800 6 la_oenb[107]
port 382 nsew signal input
rlabel metal2 s 223210 0 223266 800 6 la_oenb[108]
port 383 nsew signal input
rlabel metal2 s 224774 0 224830 800 6 la_oenb[109]
port 384 nsew signal input
rlabel metal2 s 71410 0 71466 800 6 la_oenb[10]
port 385 nsew signal input
rlabel metal2 s 226338 0 226394 800 6 la_oenb[110]
port 386 nsew signal input
rlabel metal2 s 227902 0 227958 800 6 la_oenb[111]
port 387 nsew signal input
rlabel metal2 s 229374 0 229430 800 6 la_oenb[112]
port 388 nsew signal input
rlabel metal2 s 230938 0 230994 800 6 la_oenb[113]
port 389 nsew signal input
rlabel metal2 s 232502 0 232558 800 6 la_oenb[114]
port 390 nsew signal input
rlabel metal2 s 234066 0 234122 800 6 la_oenb[115]
port 391 nsew signal input
rlabel metal2 s 235630 0 235686 800 6 la_oenb[116]
port 392 nsew signal input
rlabel metal2 s 237194 0 237250 800 6 la_oenb[117]
port 393 nsew signal input
rlabel metal2 s 238758 0 238814 800 6 la_oenb[118]
port 394 nsew signal input
rlabel metal2 s 240230 0 240286 800 6 la_oenb[119]
port 395 nsew signal input
rlabel metal2 s 72974 0 73030 800 6 la_oenb[11]
port 396 nsew signal input
rlabel metal2 s 241794 0 241850 800 6 la_oenb[120]
port 397 nsew signal input
rlabel metal2 s 243358 0 243414 800 6 la_oenb[121]
port 398 nsew signal input
rlabel metal2 s 244922 0 244978 800 6 la_oenb[122]
port 399 nsew signal input
rlabel metal2 s 246486 0 246542 800 6 la_oenb[123]
port 400 nsew signal input
rlabel metal2 s 248050 0 248106 800 6 la_oenb[124]
port 401 nsew signal input
rlabel metal2 s 249522 0 249578 800 6 la_oenb[125]
port 402 nsew signal input
rlabel metal2 s 251086 0 251142 800 6 la_oenb[126]
port 403 nsew signal input
rlabel metal2 s 252650 0 252706 800 6 la_oenb[127]
port 404 nsew signal input
rlabel metal2 s 74538 0 74594 800 6 la_oenb[12]
port 405 nsew signal input
rlabel metal2 s 76102 0 76158 800 6 la_oenb[13]
port 406 nsew signal input
rlabel metal2 s 77574 0 77630 800 6 la_oenb[14]
port 407 nsew signal input
rlabel metal2 s 79138 0 79194 800 6 la_oenb[15]
port 408 nsew signal input
rlabel metal2 s 80702 0 80758 800 6 la_oenb[16]
port 409 nsew signal input
rlabel metal2 s 82266 0 82322 800 6 la_oenb[17]
port 410 nsew signal input
rlabel metal2 s 83830 0 83886 800 6 la_oenb[18]
port 411 nsew signal input
rlabel metal2 s 85394 0 85450 800 6 la_oenb[19]
port 412 nsew signal input
rlabel metal2 s 57426 0 57482 800 6 la_oenb[1]
port 413 nsew signal input
rlabel metal2 s 86866 0 86922 800 6 la_oenb[20]
port 414 nsew signal input
rlabel metal2 s 88430 0 88486 800 6 la_oenb[21]
port 415 nsew signal input
rlabel metal2 s 89994 0 90050 800 6 la_oenb[22]
port 416 nsew signal input
rlabel metal2 s 91558 0 91614 800 6 la_oenb[23]
port 417 nsew signal input
rlabel metal2 s 93122 0 93178 800 6 la_oenb[24]
port 418 nsew signal input
rlabel metal2 s 94686 0 94742 800 6 la_oenb[25]
port 419 nsew signal input
rlabel metal2 s 96158 0 96214 800 6 la_oenb[26]
port 420 nsew signal input
rlabel metal2 s 97722 0 97778 800 6 la_oenb[27]
port 421 nsew signal input
rlabel metal2 s 99286 0 99342 800 6 la_oenb[28]
port 422 nsew signal input
rlabel metal2 s 100850 0 100906 800 6 la_oenb[29]
port 423 nsew signal input
rlabel metal2 s 58990 0 59046 800 6 la_oenb[2]
port 424 nsew signal input
rlabel metal2 s 102414 0 102470 800 6 la_oenb[30]
port 425 nsew signal input
rlabel metal2 s 103978 0 104034 800 6 la_oenb[31]
port 426 nsew signal input
rlabel metal2 s 105450 0 105506 800 6 la_oenb[32]
port 427 nsew signal input
rlabel metal2 s 107014 0 107070 800 6 la_oenb[33]
port 428 nsew signal input
rlabel metal2 s 108578 0 108634 800 6 la_oenb[34]
port 429 nsew signal input
rlabel metal2 s 110142 0 110198 800 6 la_oenb[35]
port 430 nsew signal input
rlabel metal2 s 111706 0 111762 800 6 la_oenb[36]
port 431 nsew signal input
rlabel metal2 s 113270 0 113326 800 6 la_oenb[37]
port 432 nsew signal input
rlabel metal2 s 114742 0 114798 800 6 la_oenb[38]
port 433 nsew signal input
rlabel metal2 s 116306 0 116362 800 6 la_oenb[39]
port 434 nsew signal input
rlabel metal2 s 60554 0 60610 800 6 la_oenb[3]
port 435 nsew signal input
rlabel metal2 s 117870 0 117926 800 6 la_oenb[40]
port 436 nsew signal input
rlabel metal2 s 119434 0 119490 800 6 la_oenb[41]
port 437 nsew signal input
rlabel metal2 s 120998 0 121054 800 6 la_oenb[42]
port 438 nsew signal input
rlabel metal2 s 122562 0 122618 800 6 la_oenb[43]
port 439 nsew signal input
rlabel metal2 s 124126 0 124182 800 6 la_oenb[44]
port 440 nsew signal input
rlabel metal2 s 125598 0 125654 800 6 la_oenb[45]
port 441 nsew signal input
rlabel metal2 s 127162 0 127218 800 6 la_oenb[46]
port 442 nsew signal input
rlabel metal2 s 128726 0 128782 800 6 la_oenb[47]
port 443 nsew signal input
rlabel metal2 s 130290 0 130346 800 6 la_oenb[48]
port 444 nsew signal input
rlabel metal2 s 131854 0 131910 800 6 la_oenb[49]
port 445 nsew signal input
rlabel metal2 s 62118 0 62174 800 6 la_oenb[4]
port 446 nsew signal input
rlabel metal2 s 133418 0 133474 800 6 la_oenb[50]
port 447 nsew signal input
rlabel metal2 s 134890 0 134946 800 6 la_oenb[51]
port 448 nsew signal input
rlabel metal2 s 136454 0 136510 800 6 la_oenb[52]
port 449 nsew signal input
rlabel metal2 s 138018 0 138074 800 6 la_oenb[53]
port 450 nsew signal input
rlabel metal2 s 139582 0 139638 800 6 la_oenb[54]
port 451 nsew signal input
rlabel metal2 s 141146 0 141202 800 6 la_oenb[55]
port 452 nsew signal input
rlabel metal2 s 142710 0 142766 800 6 la_oenb[56]
port 453 nsew signal input
rlabel metal2 s 144182 0 144238 800 6 la_oenb[57]
port 454 nsew signal input
rlabel metal2 s 145746 0 145802 800 6 la_oenb[58]
port 455 nsew signal input
rlabel metal2 s 147310 0 147366 800 6 la_oenb[59]
port 456 nsew signal input
rlabel metal2 s 63682 0 63738 800 6 la_oenb[5]
port 457 nsew signal input
rlabel metal2 s 148874 0 148930 800 6 la_oenb[60]
port 458 nsew signal input
rlabel metal2 s 150438 0 150494 800 6 la_oenb[61]
port 459 nsew signal input
rlabel metal2 s 152002 0 152058 800 6 la_oenb[62]
port 460 nsew signal input
rlabel metal2 s 153474 0 153530 800 6 la_oenb[63]
port 461 nsew signal input
rlabel metal2 s 155038 0 155094 800 6 la_oenb[64]
port 462 nsew signal input
rlabel metal2 s 156602 0 156658 800 6 la_oenb[65]
port 463 nsew signal input
rlabel metal2 s 158166 0 158222 800 6 la_oenb[66]
port 464 nsew signal input
rlabel metal2 s 159730 0 159786 800 6 la_oenb[67]
port 465 nsew signal input
rlabel metal2 s 161294 0 161350 800 6 la_oenb[68]
port 466 nsew signal input
rlabel metal2 s 162766 0 162822 800 6 la_oenb[69]
port 467 nsew signal input
rlabel metal2 s 65246 0 65302 800 6 la_oenb[6]
port 468 nsew signal input
rlabel metal2 s 164330 0 164386 800 6 la_oenb[70]
port 469 nsew signal input
rlabel metal2 s 165894 0 165950 800 6 la_oenb[71]
port 470 nsew signal input
rlabel metal2 s 167458 0 167514 800 6 la_oenb[72]
port 471 nsew signal input
rlabel metal2 s 169022 0 169078 800 6 la_oenb[73]
port 472 nsew signal input
rlabel metal2 s 170586 0 170642 800 6 la_oenb[74]
port 473 nsew signal input
rlabel metal2 s 172058 0 172114 800 6 la_oenb[75]
port 474 nsew signal input
rlabel metal2 s 173622 0 173678 800 6 la_oenb[76]
port 475 nsew signal input
rlabel metal2 s 175186 0 175242 800 6 la_oenb[77]
port 476 nsew signal input
rlabel metal2 s 176750 0 176806 800 6 la_oenb[78]
port 477 nsew signal input
rlabel metal2 s 178314 0 178370 800 6 la_oenb[79]
port 478 nsew signal input
rlabel metal2 s 66810 0 66866 800 6 la_oenb[7]
port 479 nsew signal input
rlabel metal2 s 179878 0 179934 800 6 la_oenb[80]
port 480 nsew signal input
rlabel metal2 s 181442 0 181498 800 6 la_oenb[81]
port 481 nsew signal input
rlabel metal2 s 182914 0 182970 800 6 la_oenb[82]
port 482 nsew signal input
rlabel metal2 s 184478 0 184534 800 6 la_oenb[83]
port 483 nsew signal input
rlabel metal2 s 186042 0 186098 800 6 la_oenb[84]
port 484 nsew signal input
rlabel metal2 s 187606 0 187662 800 6 la_oenb[85]
port 485 nsew signal input
rlabel metal2 s 189170 0 189226 800 6 la_oenb[86]
port 486 nsew signal input
rlabel metal2 s 190734 0 190790 800 6 la_oenb[87]
port 487 nsew signal input
rlabel metal2 s 192206 0 192262 800 6 la_oenb[88]
port 488 nsew signal input
rlabel metal2 s 193770 0 193826 800 6 la_oenb[89]
port 489 nsew signal input
rlabel metal2 s 68282 0 68338 800 6 la_oenb[8]
port 490 nsew signal input
rlabel metal2 s 195334 0 195390 800 6 la_oenb[90]
port 491 nsew signal input
rlabel metal2 s 196898 0 196954 800 6 la_oenb[91]
port 492 nsew signal input
rlabel metal2 s 198462 0 198518 800 6 la_oenb[92]
port 493 nsew signal input
rlabel metal2 s 200026 0 200082 800 6 la_oenb[93]
port 494 nsew signal input
rlabel metal2 s 201498 0 201554 800 6 la_oenb[94]
port 495 nsew signal input
rlabel metal2 s 203062 0 203118 800 6 la_oenb[95]
port 496 nsew signal input
rlabel metal2 s 204626 0 204682 800 6 la_oenb[96]
port 497 nsew signal input
rlabel metal2 s 206190 0 206246 800 6 la_oenb[97]
port 498 nsew signal input
rlabel metal2 s 207754 0 207810 800 6 la_oenb[98]
port 499 nsew signal input
rlabel metal2 s 209318 0 209374 800 6 la_oenb[99]
port 500 nsew signal input
rlabel metal2 s 69846 0 69902 800 6 la_oenb[9]
port 501 nsew signal input
rlabel metal4 s 4208 2128 4528 304688 6 vccd1
port 502 nsew power input
rlabel metal4 s 34928 2128 35248 304688 6 vccd1
port 502 nsew power input
rlabel metal4 s 65648 2128 65968 304688 6 vccd1
port 502 nsew power input
rlabel metal4 s 96368 2128 96688 304688 6 vccd1
port 502 nsew power input
rlabel metal4 s 127088 2128 127408 304688 6 vccd1
port 502 nsew power input
rlabel metal4 s 157808 2128 158128 304688 6 vccd1
port 502 nsew power input
rlabel metal4 s 188528 2128 188848 304688 6 vccd1
port 502 nsew power input
rlabel metal4 s 219248 2128 219568 304688 6 vccd1
port 502 nsew power input
rlabel metal4 s 249968 2128 250288 304688 6 vccd1
port 502 nsew power input
rlabel metal4 s 19568 2128 19888 304688 6 vssd1
port 503 nsew ground input
rlabel metal4 s 50288 2128 50608 304688 6 vssd1
port 503 nsew ground input
rlabel metal4 s 81008 2128 81328 304688 6 vssd1
port 503 nsew ground input
rlabel metal4 s 111728 2128 112048 304688 6 vssd1
port 503 nsew ground input
rlabel metal4 s 142448 2128 142768 304688 6 vssd1
port 503 nsew ground input
rlabel metal4 s 173168 2128 173488 304688 6 vssd1
port 503 nsew ground input
rlabel metal4 s 203888 2128 204208 304688 6 vssd1
port 503 nsew ground input
rlabel metal4 s 234608 2128 234928 304688 6 vssd1
port 503 nsew ground input
rlabel metal2 s 202 0 258 800 6 wb_clk_i
port 504 nsew signal input
rlabel metal2 s 662 0 718 800 6 wb_rst_i
port 505 nsew signal input
rlabel metal2 s 1214 0 1270 800 6 wbs_ack_o
port 506 nsew signal output
rlabel metal2 s 3238 0 3294 800 6 wbs_adr_i[0]
port 507 nsew signal input
rlabel metal2 s 20810 0 20866 800 6 wbs_adr_i[10]
port 508 nsew signal input
rlabel metal2 s 22374 0 22430 800 6 wbs_adr_i[11]
port 509 nsew signal input
rlabel metal2 s 23938 0 23994 800 6 wbs_adr_i[12]
port 510 nsew signal input
rlabel metal2 s 25502 0 25558 800 6 wbs_adr_i[13]
port 511 nsew signal input
rlabel metal2 s 26974 0 27030 800 6 wbs_adr_i[14]
port 512 nsew signal input
rlabel metal2 s 28538 0 28594 800 6 wbs_adr_i[15]
port 513 nsew signal input
rlabel metal2 s 30102 0 30158 800 6 wbs_adr_i[16]
port 514 nsew signal input
rlabel metal2 s 31666 0 31722 800 6 wbs_adr_i[17]
port 515 nsew signal input
rlabel metal2 s 33230 0 33286 800 6 wbs_adr_i[18]
port 516 nsew signal input
rlabel metal2 s 34794 0 34850 800 6 wbs_adr_i[19]
port 517 nsew signal input
rlabel metal2 s 5354 0 5410 800 6 wbs_adr_i[1]
port 518 nsew signal input
rlabel metal2 s 36266 0 36322 800 6 wbs_adr_i[20]
port 519 nsew signal input
rlabel metal2 s 37830 0 37886 800 6 wbs_adr_i[21]
port 520 nsew signal input
rlabel metal2 s 39394 0 39450 800 6 wbs_adr_i[22]
port 521 nsew signal input
rlabel metal2 s 40958 0 41014 800 6 wbs_adr_i[23]
port 522 nsew signal input
rlabel metal2 s 42522 0 42578 800 6 wbs_adr_i[24]
port 523 nsew signal input
rlabel metal2 s 44086 0 44142 800 6 wbs_adr_i[25]
port 524 nsew signal input
rlabel metal2 s 45558 0 45614 800 6 wbs_adr_i[26]
port 525 nsew signal input
rlabel metal2 s 47122 0 47178 800 6 wbs_adr_i[27]
port 526 nsew signal input
rlabel metal2 s 48686 0 48742 800 6 wbs_adr_i[28]
port 527 nsew signal input
rlabel metal2 s 50250 0 50306 800 6 wbs_adr_i[29]
port 528 nsew signal input
rlabel metal2 s 7378 0 7434 800 6 wbs_adr_i[2]
port 529 nsew signal input
rlabel metal2 s 51814 0 51870 800 6 wbs_adr_i[30]
port 530 nsew signal input
rlabel metal2 s 53378 0 53434 800 6 wbs_adr_i[31]
port 531 nsew signal input
rlabel metal2 s 9494 0 9550 800 6 wbs_adr_i[3]
port 532 nsew signal input
rlabel metal2 s 11518 0 11574 800 6 wbs_adr_i[4]
port 533 nsew signal input
rlabel metal2 s 13082 0 13138 800 6 wbs_adr_i[5]
port 534 nsew signal input
rlabel metal2 s 14646 0 14702 800 6 wbs_adr_i[6]
port 535 nsew signal input
rlabel metal2 s 16118 0 16174 800 6 wbs_adr_i[7]
port 536 nsew signal input
rlabel metal2 s 17682 0 17738 800 6 wbs_adr_i[8]
port 537 nsew signal input
rlabel metal2 s 19246 0 19302 800 6 wbs_adr_i[9]
port 538 nsew signal input
rlabel metal2 s 1674 0 1730 800 6 wbs_cyc_i
port 539 nsew signal input
rlabel metal2 s 3790 0 3846 800 6 wbs_dat_i[0]
port 540 nsew signal input
rlabel metal2 s 21362 0 21418 800 6 wbs_dat_i[10]
port 541 nsew signal input
rlabel metal2 s 22834 0 22890 800 6 wbs_dat_i[11]
port 542 nsew signal input
rlabel metal2 s 24398 0 24454 800 6 wbs_dat_i[12]
port 543 nsew signal input
rlabel metal2 s 25962 0 26018 800 6 wbs_dat_i[13]
port 544 nsew signal input
rlabel metal2 s 27526 0 27582 800 6 wbs_dat_i[14]
port 545 nsew signal input
rlabel metal2 s 29090 0 29146 800 6 wbs_dat_i[15]
port 546 nsew signal input
rlabel metal2 s 30654 0 30710 800 6 wbs_dat_i[16]
port 547 nsew signal input
rlabel metal2 s 32126 0 32182 800 6 wbs_dat_i[17]
port 548 nsew signal input
rlabel metal2 s 33690 0 33746 800 6 wbs_dat_i[18]
port 549 nsew signal input
rlabel metal2 s 35254 0 35310 800 6 wbs_dat_i[19]
port 550 nsew signal input
rlabel metal2 s 5814 0 5870 800 6 wbs_dat_i[1]
port 551 nsew signal input
rlabel metal2 s 36818 0 36874 800 6 wbs_dat_i[20]
port 552 nsew signal input
rlabel metal2 s 38382 0 38438 800 6 wbs_dat_i[21]
port 553 nsew signal input
rlabel metal2 s 39946 0 40002 800 6 wbs_dat_i[22]
port 554 nsew signal input
rlabel metal2 s 41510 0 41566 800 6 wbs_dat_i[23]
port 555 nsew signal input
rlabel metal2 s 42982 0 43038 800 6 wbs_dat_i[24]
port 556 nsew signal input
rlabel metal2 s 44546 0 44602 800 6 wbs_dat_i[25]
port 557 nsew signal input
rlabel metal2 s 46110 0 46166 800 6 wbs_dat_i[26]
port 558 nsew signal input
rlabel metal2 s 47674 0 47730 800 6 wbs_dat_i[27]
port 559 nsew signal input
rlabel metal2 s 49238 0 49294 800 6 wbs_dat_i[28]
port 560 nsew signal input
rlabel metal2 s 50802 0 50858 800 6 wbs_dat_i[29]
port 561 nsew signal input
rlabel metal2 s 7930 0 7986 800 6 wbs_dat_i[2]
port 562 nsew signal input
rlabel metal2 s 52274 0 52330 800 6 wbs_dat_i[30]
port 563 nsew signal input
rlabel metal2 s 53838 0 53894 800 6 wbs_dat_i[31]
port 564 nsew signal input
rlabel metal2 s 9954 0 10010 800 6 wbs_dat_i[3]
port 565 nsew signal input
rlabel metal2 s 12070 0 12126 800 6 wbs_dat_i[4]
port 566 nsew signal input
rlabel metal2 s 13542 0 13598 800 6 wbs_dat_i[5]
port 567 nsew signal input
rlabel metal2 s 15106 0 15162 800 6 wbs_dat_i[6]
port 568 nsew signal input
rlabel metal2 s 16670 0 16726 800 6 wbs_dat_i[7]
port 569 nsew signal input
rlabel metal2 s 18234 0 18290 800 6 wbs_dat_i[8]
port 570 nsew signal input
rlabel metal2 s 19798 0 19854 800 6 wbs_dat_i[9]
port 571 nsew signal input
rlabel metal2 s 4250 0 4306 800 6 wbs_dat_o[0]
port 572 nsew signal output
rlabel metal2 s 21822 0 21878 800 6 wbs_dat_o[10]
port 573 nsew signal output
rlabel metal2 s 23386 0 23442 800 6 wbs_dat_o[11]
port 574 nsew signal output
rlabel metal2 s 24950 0 25006 800 6 wbs_dat_o[12]
port 575 nsew signal output
rlabel metal2 s 26514 0 26570 800 6 wbs_dat_o[13]
port 576 nsew signal output
rlabel metal2 s 28078 0 28134 800 6 wbs_dat_o[14]
port 577 nsew signal output
rlabel metal2 s 29550 0 29606 800 6 wbs_dat_o[15]
port 578 nsew signal output
rlabel metal2 s 31114 0 31170 800 6 wbs_dat_o[16]
port 579 nsew signal output
rlabel metal2 s 32678 0 32734 800 6 wbs_dat_o[17]
port 580 nsew signal output
rlabel metal2 s 34242 0 34298 800 6 wbs_dat_o[18]
port 581 nsew signal output
rlabel metal2 s 35806 0 35862 800 6 wbs_dat_o[19]
port 582 nsew signal output
rlabel metal2 s 6366 0 6422 800 6 wbs_dat_o[1]
port 583 nsew signal output
rlabel metal2 s 37370 0 37426 800 6 wbs_dat_o[20]
port 584 nsew signal output
rlabel metal2 s 38842 0 38898 800 6 wbs_dat_o[21]
port 585 nsew signal output
rlabel metal2 s 40406 0 40462 800 6 wbs_dat_o[22]
port 586 nsew signal output
rlabel metal2 s 41970 0 42026 800 6 wbs_dat_o[23]
port 587 nsew signal output
rlabel metal2 s 43534 0 43590 800 6 wbs_dat_o[24]
port 588 nsew signal output
rlabel metal2 s 45098 0 45154 800 6 wbs_dat_o[25]
port 589 nsew signal output
rlabel metal2 s 46662 0 46718 800 6 wbs_dat_o[26]
port 590 nsew signal output
rlabel metal2 s 48134 0 48190 800 6 wbs_dat_o[27]
port 591 nsew signal output
rlabel metal2 s 49698 0 49754 800 6 wbs_dat_o[28]
port 592 nsew signal output
rlabel metal2 s 51262 0 51318 800 6 wbs_dat_o[29]
port 593 nsew signal output
rlabel metal2 s 8390 0 8446 800 6 wbs_dat_o[2]
port 594 nsew signal output
rlabel metal2 s 52826 0 52882 800 6 wbs_dat_o[30]
port 595 nsew signal output
rlabel metal2 s 54390 0 54446 800 6 wbs_dat_o[31]
port 596 nsew signal output
rlabel metal2 s 10506 0 10562 800 6 wbs_dat_o[3]
port 597 nsew signal output
rlabel metal2 s 12530 0 12586 800 6 wbs_dat_o[4]
port 598 nsew signal output
rlabel metal2 s 14094 0 14150 800 6 wbs_dat_o[5]
port 599 nsew signal output
rlabel metal2 s 15658 0 15714 800 6 wbs_dat_o[6]
port 600 nsew signal output
rlabel metal2 s 17222 0 17278 800 6 wbs_dat_o[7]
port 601 nsew signal output
rlabel metal2 s 18786 0 18842 800 6 wbs_dat_o[8]
port 602 nsew signal output
rlabel metal2 s 20258 0 20314 800 6 wbs_dat_o[9]
port 603 nsew signal output
rlabel metal2 s 4802 0 4858 800 6 wbs_sel_i[0]
port 604 nsew signal input
rlabel metal2 s 6826 0 6882 800 6 wbs_sel_i[1]
port 605 nsew signal input
rlabel metal2 s 8942 0 8998 800 6 wbs_sel_i[2]
port 606 nsew signal input
rlabel metal2 s 10966 0 11022 800 6 wbs_sel_i[3]
port 607 nsew signal input
rlabel metal2 s 2226 0 2282 800 6 wbs_stb_i
port 608 nsew signal input
rlabel metal2 s 2778 0 2834 800 6 wbs_we_i
port 609 nsew signal input
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 254531 307139
string LEFview TRUE
string GDS_FILE /project/openlane/user_project/runs/user_project/results/magic/user_project.gds
string GDS_END 249570672
string GDS_START 1071792
<< end >>

