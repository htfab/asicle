magic
tech sky130A
magscale 1 2
timestamp 1647846298
<< locali >>
rect 205097 506651 205131 507569
rect 218529 506719 218563 507637
rect 237389 507127 237423 509201
rect 349571 507229 349905 507263
rect 349663 507161 349813 507195
rect 349571 507093 349905 507127
rect 356713 506991 356747 508453
rect 358921 506855 358955 508453
rect 363337 506923 363371 508453
rect 370053 506787 370087 508317
rect 383485 506583 383519 508181
rect 396549 506515 396583 507977
rect 400079 198645 400171 198679
rect 201509 198441 201693 198475
rect 201509 198407 201543 198441
rect 394893 197591 394927 197829
rect 397101 197523 397135 197761
rect 400137 197387 400171 198645
rect 407773 197795 407807 197897
rect 420193 197523 420227 198509
rect 428657 197455 428691 197557
rect 327549 4743 327583 5049
rect 416513 5049 416973 5083
rect 416513 4947 416547 5049
rect 416823 4981 417065 5015
rect 368891 4165 369133 4199
rect 175933 3961 176117 3995
rect 175933 3927 175967 3961
rect 164801 3451 164835 3689
rect 240425 3383 240459 3485
rect 253213 3451 253247 3961
rect 258181 3859 258215 4029
rect 312461 3927 312495 4097
rect 258123 3825 258215 3859
rect 314025 3655 314059 3825
rect 317521 3519 317555 3689
rect 320833 3315 320867 3689
rect 360025 3179 360059 3553
rect 368949 3315 368983 4097
<< viali >>
rect 237389 509201 237423 509235
rect 218529 507637 218563 507671
rect 205097 507569 205131 507603
rect 356713 508453 356747 508487
rect 349537 507229 349571 507263
rect 349905 507229 349939 507263
rect 349629 507161 349663 507195
rect 349813 507161 349847 507195
rect 237389 507093 237423 507127
rect 349537 507093 349571 507127
rect 349905 507093 349939 507127
rect 356713 506957 356747 506991
rect 358921 508453 358955 508487
rect 363337 508453 363371 508487
rect 363337 506889 363371 506923
rect 370053 508317 370087 508351
rect 358921 506821 358955 506855
rect 370053 506753 370087 506787
rect 383485 508181 383519 508215
rect 218529 506685 218563 506719
rect 205097 506617 205131 506651
rect 383485 506549 383519 506583
rect 396549 507977 396583 508011
rect 396549 506481 396583 506515
rect 400045 198645 400079 198679
rect 201693 198441 201727 198475
rect 201509 198373 201543 198407
rect 394893 197829 394927 197863
rect 394893 197557 394927 197591
rect 397101 197761 397135 197795
rect 397101 197489 397135 197523
rect 420193 198509 420227 198543
rect 407773 197897 407807 197931
rect 407773 197761 407807 197795
rect 420193 197489 420227 197523
rect 428657 197557 428691 197591
rect 428657 197421 428691 197455
rect 400137 197353 400171 197387
rect 327549 5049 327583 5083
rect 416973 5049 417007 5083
rect 416789 4981 416823 5015
rect 417065 4981 417099 5015
rect 416513 4913 416547 4947
rect 327549 4709 327583 4743
rect 368857 4165 368891 4199
rect 369133 4165 369167 4199
rect 312461 4097 312495 4131
rect 258181 4029 258215 4063
rect 176117 3961 176151 3995
rect 253213 3961 253247 3995
rect 175933 3893 175967 3927
rect 164801 3689 164835 3723
rect 164801 3417 164835 3451
rect 240425 3485 240459 3519
rect 312461 3893 312495 3927
rect 368949 4097 368983 4131
rect 258089 3825 258123 3859
rect 314025 3825 314059 3859
rect 314025 3621 314059 3655
rect 317521 3689 317555 3723
rect 317521 3485 317555 3519
rect 320833 3689 320867 3723
rect 253213 3417 253247 3451
rect 240425 3349 240459 3383
rect 320833 3281 320867 3315
rect 360025 3553 360059 3587
rect 368949 3281 368983 3315
rect 360025 3145 360059 3179
<< metal1 >>
rect 137830 700952 137836 701004
rect 137888 700992 137894 701004
rect 309134 700992 309140 701004
rect 137888 700964 309140 700992
rect 137888 700952 137894 700964
rect 309134 700952 309140 700964
rect 309192 700952 309198 701004
rect 277302 700884 277308 700936
rect 277360 700924 277366 700936
rect 462314 700924 462320 700936
rect 277360 700896 462320 700924
rect 277360 700884 277366 700896
rect 462314 700884 462320 700896
rect 462372 700884 462378 700936
rect 278682 700816 278688 700868
rect 278740 700856 278746 700868
rect 478506 700856 478512 700868
rect 278740 700828 478512 700856
rect 278740 700816 278746 700828
rect 478506 700816 478512 700828
rect 478564 700816 478570 700868
rect 105446 700748 105452 700800
rect 105504 700788 105510 700800
rect 313274 700788 313280 700800
rect 105504 700760 313280 700788
rect 105504 700748 105510 700760
rect 313274 700748 313280 700760
rect 313332 700748 313338 700800
rect 89162 700680 89168 700732
rect 89220 700720 89226 700732
rect 317414 700720 317420 700732
rect 89220 700692 317420 700720
rect 89220 700680 89226 700692
rect 317414 700680 317420 700692
rect 317472 700680 317478 700732
rect 72970 700612 72976 700664
rect 73028 700652 73034 700664
rect 316034 700652 316040 700664
rect 73028 700624 316040 700652
rect 73028 700612 73034 700624
rect 316034 700612 316040 700624
rect 316092 700612 316098 700664
rect 270402 700544 270408 700596
rect 270460 700584 270466 700596
rect 527174 700584 527180 700596
rect 270460 700556 527180 700584
rect 270460 700544 270466 700556
rect 527174 700544 527180 700556
rect 527232 700544 527238 700596
rect 271782 700476 271788 700528
rect 271840 700516 271846 700528
rect 543458 700516 543464 700528
rect 271840 700488 543464 700516
rect 271840 700476 271846 700488
rect 543458 700476 543464 700488
rect 543516 700476 543522 700528
rect 40494 700408 40500 700460
rect 40552 700448 40558 700460
rect 320174 700448 320180 700460
rect 40552 700420 320180 700448
rect 40552 700408 40558 700420
rect 320174 700408 320180 700420
rect 320232 700408 320238 700460
rect 24302 700340 24308 700392
rect 24360 700380 24366 700392
rect 324314 700380 324320 700392
rect 24360 700352 324320 700380
rect 24360 700340 24366 700352
rect 324314 700340 324320 700352
rect 324372 700340 324378 700392
rect 8110 700272 8116 700324
rect 8168 700312 8174 700324
rect 322934 700312 322940 700324
rect 8168 700284 322940 700312
rect 8168 700272 8174 700284
rect 322934 700272 322940 700284
rect 322992 700272 322998 700324
rect 154114 700204 154120 700256
rect 154172 700244 154178 700256
rect 311894 700244 311900 700256
rect 154172 700216 311900 700244
rect 154172 700204 154178 700216
rect 311894 700204 311900 700216
rect 311952 700204 311958 700256
rect 285582 700136 285588 700188
rect 285640 700176 285646 700188
rect 413646 700176 413652 700188
rect 285640 700148 413652 700176
rect 285640 700136 285646 700148
rect 413646 700136 413652 700148
rect 413704 700136 413710 700188
rect 202782 700068 202788 700120
rect 202840 700108 202846 700120
rect 302234 700108 302240 700120
rect 202840 700080 302240 700108
rect 202840 700068 202846 700080
rect 302234 700068 302240 700080
rect 302292 700068 302298 700120
rect 302878 700068 302884 700120
rect 302936 700108 302942 700120
rect 429838 700108 429844 700120
rect 302936 700080 429844 700108
rect 302936 700068 302942 700080
rect 429838 700068 429844 700080
rect 429896 700068 429902 700120
rect 284202 700000 284208 700052
rect 284260 700040 284266 700052
rect 397454 700040 397460 700052
rect 284260 700012 397460 700040
rect 284260 700000 284266 700012
rect 397454 700000 397460 700012
rect 397512 700000 397518 700052
rect 292482 699932 292488 699984
rect 292540 699972 292546 699984
rect 348786 699972 348792 699984
rect 292540 699944 348792 699972
rect 292540 699932 292546 699944
rect 348786 699932 348792 699944
rect 348844 699932 348850 699984
rect 289722 699864 289728 699916
rect 289780 699904 289786 699916
rect 332502 699904 332508 699916
rect 289780 699876 332508 699904
rect 289780 699864 289786 699876
rect 332502 699864 332508 699876
rect 332560 699864 332566 699916
rect 267642 699796 267648 699848
rect 267700 699836 267706 699848
rect 295334 699836 295340 699848
rect 267700 699808 295340 699836
rect 267700 699796 267706 699808
rect 295334 699796 295340 699808
rect 295392 699796 295398 699848
rect 283834 699728 283840 699780
rect 283892 699768 283898 699780
rect 298094 699768 298100 699780
rect 283892 699740 298100 699768
rect 283892 699728 283898 699740
rect 298094 699728 298100 699740
rect 298152 699728 298158 699780
rect 170306 699660 170312 699712
rect 170364 699700 170370 699712
rect 171042 699700 171048 699712
rect 170364 699672 171048 699700
rect 170364 699660 170370 699672
rect 171042 699660 171048 699672
rect 171100 699660 171106 699712
rect 235166 699660 235172 699712
rect 235224 699700 235230 699712
rect 235902 699700 235908 699712
rect 235224 699672 235908 699700
rect 235224 699660 235230 699672
rect 235902 699660 235908 699672
rect 235960 699660 235966 699712
rect 263502 696940 263508 696992
rect 263560 696980 263566 696992
rect 580166 696980 580172 696992
rect 263560 696952 580172 696980
rect 263560 696940 263566 696952
rect 580166 696940 580172 696952
rect 580224 696940 580230 696992
rect 266262 683204 266268 683256
rect 266320 683244 266326 683256
rect 580166 683244 580172 683256
rect 266320 683216 580172 683244
rect 266320 683204 266326 683216
rect 580166 683204 580172 683216
rect 580224 683204 580230 683256
rect 3418 683136 3424 683188
rect 3476 683176 3482 683188
rect 327074 683176 327080 683188
rect 3476 683148 327080 683176
rect 3476 683136 3482 683148
rect 327074 683136 327080 683148
rect 327132 683136 327138 683188
rect 260742 670760 260748 670812
rect 260800 670800 260806 670812
rect 580166 670800 580172 670812
rect 260800 670772 580172 670800
rect 260800 670760 260806 670772
rect 580166 670760 580172 670772
rect 580224 670760 580230 670812
rect 3510 670692 3516 670744
rect 3568 670732 3574 670744
rect 331214 670732 331220 670744
rect 3568 670704 331220 670732
rect 3568 670692 3574 670704
rect 331214 670692 331220 670704
rect 331272 670692 331278 670744
rect 3418 656888 3424 656940
rect 3476 656928 3482 656940
rect 329834 656928 329840 656940
rect 3476 656900 329840 656928
rect 3476 656888 3482 656900
rect 329834 656888 329840 656900
rect 329892 656888 329898 656940
rect 256602 643084 256608 643136
rect 256660 643124 256666 643136
rect 580166 643124 580172 643136
rect 256660 643096 580172 643124
rect 256660 643084 256666 643096
rect 580166 643084 580172 643096
rect 580224 643084 580230 643136
rect 3418 632068 3424 632120
rect 3476 632108 3482 632120
rect 333974 632108 333980 632120
rect 3476 632080 333980 632108
rect 3476 632068 3482 632080
rect 333974 632068 333980 632080
rect 334032 632068 334038 632120
rect 259362 630640 259368 630692
rect 259420 630680 259426 630692
rect 580166 630680 580172 630692
rect 259420 630652 580172 630680
rect 259420 630640 259426 630652
rect 580166 630640 580172 630652
rect 580224 630640 580230 630692
rect 3142 618264 3148 618316
rect 3200 618304 3206 618316
rect 338114 618304 338120 618316
rect 3200 618276 338120 618304
rect 3200 618264 3206 618276
rect 338114 618264 338120 618276
rect 338172 618264 338178 618316
rect 255222 616836 255228 616888
rect 255280 616876 255286 616888
rect 580166 616876 580172 616888
rect 255280 616848 580172 616876
rect 255280 616836 255286 616848
rect 580166 616836 580172 616848
rect 580224 616836 580230 616888
rect 3234 605820 3240 605872
rect 3292 605860 3298 605872
rect 335354 605860 335360 605872
rect 3292 605832 335360 605860
rect 3292 605820 3298 605832
rect 335354 605820 335360 605832
rect 335412 605820 335418 605872
rect 249702 590656 249708 590708
rect 249760 590696 249766 590708
rect 579798 590696 579804 590708
rect 249760 590668 579804 590696
rect 249760 590656 249766 590668
rect 579798 590656 579804 590668
rect 579856 590656 579862 590708
rect 3326 579640 3332 579692
rect 3384 579680 3390 579692
rect 340874 579680 340880 579692
rect 3384 579652 340880 579680
rect 3384 579640 3390 579652
rect 340874 579640 340880 579652
rect 340932 579640 340938 579692
rect 252462 576852 252468 576904
rect 252520 576892 252526 576904
rect 580166 576892 580172 576904
rect 252520 576864 580172 576892
rect 252520 576852 252526 576864
rect 580166 576852 580172 576864
rect 580224 576852 580230 576904
rect 3418 565836 3424 565888
rect 3476 565876 3482 565888
rect 345014 565876 345020 565888
rect 3476 565848 345020 565876
rect 3476 565836 3482 565848
rect 345014 565836 345020 565848
rect 345072 565836 345078 565888
rect 248322 563048 248328 563100
rect 248380 563088 248386 563100
rect 579798 563088 579804 563100
rect 248380 563060 579804 563088
rect 248380 563048 248386 563060
rect 579798 563048 579804 563060
rect 579856 563048 579862 563100
rect 3418 553392 3424 553444
rect 3476 553432 3482 553444
rect 342254 553432 342260 553444
rect 3476 553404 342260 553432
rect 3476 553392 3482 553404
rect 342254 553392 342260 553404
rect 342312 553392 342318 553444
rect 242802 536800 242808 536852
rect 242860 536840 242866 536852
rect 580166 536840 580172 536852
rect 242860 536812 580172 536840
rect 242860 536800 242866 536812
rect 580166 536800 580172 536812
rect 580224 536800 580230 536852
rect 3418 527144 3424 527196
rect 3476 527184 3482 527196
rect 347774 527184 347780 527196
rect 3476 527156 347780 527184
rect 3476 527144 3482 527156
rect 347774 527144 347780 527156
rect 347832 527144 347838 527196
rect 245562 524424 245568 524476
rect 245620 524464 245626 524476
rect 580166 524464 580172 524476
rect 245620 524436 580172 524464
rect 245620 524424 245626 524436
rect 580166 524424 580172 524436
rect 580224 524424 580230 524476
rect 3418 514768 3424 514820
rect 3476 514808 3482 514820
rect 351914 514808 351920 514820
rect 3476 514780 351920 514808
rect 3476 514768 3482 514780
rect 351914 514768 351920 514780
rect 351972 514768 351978 514820
rect 294138 511708 294144 511760
rect 294196 511748 294202 511760
rect 299474 511748 299480 511760
rect 294196 511720 299480 511748
rect 294196 511708 294202 511720
rect 299474 511708 299480 511720
rect 299532 511708 299538 511760
rect 280706 511640 280712 511692
rect 280764 511680 280770 511692
rect 302878 511680 302884 511692
rect 280764 511652 302884 511680
rect 280764 511640 280770 511652
rect 302878 511640 302884 511652
rect 302936 511640 302942 511692
rect 235902 511572 235908 511624
rect 235960 511612 235966 511624
rect 300854 511612 300860 511624
rect 235960 511584 300860 511612
rect 235960 511572 235966 511584
rect 300854 511572 300860 511584
rect 300912 511572 300918 511624
rect 287422 511504 287428 511556
rect 287480 511544 287486 511556
rect 364334 511544 364340 511556
rect 287480 511516 364340 511544
rect 287480 511504 287486 511516
rect 364334 511504 364340 511516
rect 364392 511504 364398 511556
rect 219342 511436 219348 511488
rect 219400 511476 219406 511488
rect 305270 511476 305276 511488
rect 219400 511448 305276 511476
rect 219400 511436 219406 511448
rect 305270 511436 305276 511448
rect 305328 511436 305334 511488
rect 171042 511368 171048 511420
rect 171100 511408 171106 511420
rect 307570 511408 307576 511420
rect 171100 511380 307576 511408
rect 171100 511368 171106 511380
rect 307570 511368 307576 511380
rect 307628 511368 307634 511420
rect 274082 511300 274088 511352
rect 274140 511340 274146 511352
rect 494054 511340 494060 511352
rect 274140 511312 494060 511340
rect 274140 511300 274146 511312
rect 494054 511300 494060 511312
rect 494112 511300 494118 511352
rect 267366 511232 267372 511284
rect 267424 511272 267430 511284
rect 558914 511272 558920 511284
rect 267424 511244 558920 511272
rect 267424 511232 267430 511244
rect 558914 511232 558920 511244
rect 558972 511232 558978 511284
rect 240502 510620 240508 510672
rect 240560 510660 240566 510672
rect 580166 510660 580172 510672
rect 240560 510632 580172 510660
rect 240560 510620 240566 510632
rect 580166 510620 580172 510632
rect 580224 510620 580230 510672
rect 198090 510552 198096 510604
rect 198148 510592 198154 510604
rect 237374 510592 237380 510604
rect 198148 510564 237380 510592
rect 198148 510552 198154 510564
rect 237374 510552 237380 510564
rect 237432 510552 237438 510604
rect 238294 510552 238300 510604
rect 238352 510592 238358 510604
rect 431310 510592 431316 510604
rect 238352 510564 431316 510592
rect 238352 510552 238358 510564
rect 431310 510552 431316 510564
rect 431368 510552 431374 510604
rect 231578 510484 231584 510536
rect 231636 510524 231642 510536
rect 431218 510524 431224 510536
rect 231636 510496 431224 510524
rect 231636 510484 231642 510496
rect 431218 510484 431224 510496
rect 431276 510484 431282 510536
rect 229370 510416 229376 510468
rect 229428 510456 229434 510468
rect 430114 510456 430120 510468
rect 229428 510428 430120 510456
rect 229428 510416 229434 510428
rect 430114 510416 430120 510428
rect 430172 510416 430178 510468
rect 175826 510348 175832 510400
rect 175884 510388 175890 510400
rect 424318 510388 424324 510400
rect 175884 510360 424324 510388
rect 175884 510348 175890 510360
rect 424318 510348 424324 510360
rect 424376 510348 424382 510400
rect 215938 510280 215944 510332
rect 215996 510320 216002 510332
rect 478138 510320 478144 510332
rect 215996 510292 478144 510320
rect 215996 510280 216002 510292
rect 478138 510280 478144 510292
rect 478196 510280 478202 510332
rect 224954 510212 224960 510264
rect 225012 510252 225018 510264
rect 496078 510252 496084 510264
rect 225012 510224 496084 510252
rect 225012 510212 225018 510224
rect 496078 510212 496084 510224
rect 496136 510212 496142 510264
rect 100110 510144 100116 510196
rect 100168 510184 100174 510196
rect 399110 510184 399116 510196
rect 100168 510156 399116 510184
rect 100168 510144 100174 510156
rect 399110 510144 399116 510156
rect 399168 510144 399174 510196
rect 101490 510076 101496 510128
rect 101548 510116 101554 510128
rect 405826 510116 405832 510128
rect 101548 510088 405832 510116
rect 101548 510076 101554 510088
rect 405826 510076 405832 510088
rect 405884 510076 405890 510128
rect 100018 510008 100024 510060
rect 100076 510048 100082 510060
rect 412450 510048 412456 510060
rect 100076 510020 412456 510048
rect 100076 510008 100082 510020
rect 412450 510008 412456 510020
rect 412508 510008 412514 510060
rect 101398 509940 101404 509992
rect 101456 509980 101462 509992
rect 419166 509980 419172 509992
rect 101456 509952 419172 509980
rect 101456 509940 101462 509952
rect 419166 509940 419172 509952
rect 419224 509940 419230 509992
rect 82078 509872 82084 509924
rect 82136 509912 82142 509924
rect 410242 509912 410248 509924
rect 82136 509884 410248 509912
rect 82136 509872 82142 509884
rect 410242 509872 410248 509884
rect 410300 509872 410306 509924
rect 64138 509804 64144 509856
rect 64196 509844 64202 509856
rect 403526 509844 403532 509856
rect 64196 509816 403532 509844
rect 64196 509804 64202 509816
rect 403526 509804 403532 509816
rect 403584 509804 403590 509856
rect 222654 509736 222660 509788
rect 222712 509776 222718 509788
rect 562318 509776 562324 509788
rect 222712 509748 562324 509776
rect 222712 509736 222718 509748
rect 562318 509736 562324 509748
rect 562376 509736 562382 509788
rect 4982 509668 4988 509720
rect 5040 509708 5046 509720
rect 365622 509708 365628 509720
rect 5040 509680 365628 509708
rect 5040 509668 5046 509680
rect 365622 509668 365628 509680
rect 365680 509668 365686 509720
rect 14642 509600 14648 509652
rect 14700 509640 14706 509652
rect 376754 509640 376760 509652
rect 14700 509612 376760 509640
rect 14700 509600 14706 509612
rect 376754 509600 376760 509612
rect 376812 509600 376818 509652
rect 4890 509532 4896 509584
rect 4948 509572 4954 509584
rect 372338 509572 372344 509584
rect 4948 509544 372344 509572
rect 4948 509532 4954 509544
rect 372338 509532 372344 509544
rect 372396 509532 372402 509584
rect 11698 509464 11704 509516
rect 11756 509504 11762 509516
rect 378962 509504 378968 509516
rect 11756 509476 378968 509504
rect 11756 509464 11762 509476
rect 378962 509464 378968 509476
rect 379020 509464 379026 509516
rect 14550 509396 14556 509448
rect 14608 509436 14614 509448
rect 385678 509436 385684 509448
rect 14608 509408 385684 509436
rect 14608 509396 14614 509408
rect 385678 509396 385684 509408
rect 385736 509396 385742 509448
rect 14458 509328 14464 509380
rect 14516 509368 14522 509380
rect 392394 509368 392400 509380
rect 14516 509340 392400 509368
rect 14516 509328 14522 509340
rect 392394 509328 392400 509340
rect 392452 509328 392458 509380
rect 4798 509260 4804 509312
rect 4856 509300 4862 509312
rect 390186 509300 390192 509312
rect 4856 509272 390192 509300
rect 4856 509260 4862 509272
rect 390186 509260 390192 509272
rect 390244 509260 390250 509312
rect 237374 509232 237380 509244
rect 237335 509204 237380 509232
rect 237374 509192 237380 509204
rect 237432 509192 237438 509244
rect 233878 509124 233884 509176
rect 233936 509164 233942 509176
rect 421926 509164 421932 509176
rect 233936 509136 421932 509164
rect 233936 509124 233942 509136
rect 421926 509124 421932 509136
rect 421984 509124 421990 509176
rect 213730 509056 213736 509108
rect 213788 509096 213794 509108
rect 425882 509096 425888 509108
rect 213788 509068 425888 509096
rect 213788 509056 213794 509068
rect 425882 509056 425888 509068
rect 425940 509056 425946 509108
rect 207014 508988 207020 509040
rect 207072 509028 207078 509040
rect 424502 509028 424508 509040
rect 207072 509000 424508 509028
rect 207072 508988 207078 509000
rect 424502 508988 424508 509000
rect 424560 508988 424566 509040
rect 200390 508920 200396 508972
rect 200448 508960 200454 508972
rect 422938 508960 422944 508972
rect 200448 508932 422944 508960
rect 200448 508920 200454 508932
rect 422938 508920 422944 508932
rect 422996 508920 423002 508972
rect 193674 508852 193680 508904
rect 193732 508892 193738 508904
rect 424410 508892 424416 508904
rect 193732 508864 424416 508892
rect 193732 508852 193738 508864
rect 424410 508852 424416 508864
rect 424468 508852 424474 508904
rect 186958 508784 186964 508836
rect 187016 508824 187022 508836
rect 421834 508824 421840 508836
rect 187016 508796 421840 508824
rect 187016 508784 187022 508796
rect 421834 508784 421840 508796
rect 421892 508784 421898 508836
rect 180242 508716 180248 508768
rect 180300 508756 180306 508768
rect 421742 508756 421748 508768
rect 180300 508728 421748 508756
rect 180300 508716 180306 508728
rect 421742 508716 421748 508728
rect 421800 508716 421806 508768
rect 173526 508648 173532 508700
rect 173584 508688 173590 508700
rect 421650 508688 421656 508700
rect 173584 508660 421656 508688
rect 173584 508648 173590 508660
rect 421650 508648 421656 508660
rect 421708 508648 421714 508700
rect 169110 508580 169116 508632
rect 169168 508620 169174 508632
rect 508498 508620 508504 508632
rect 169168 508592 508504 508620
rect 169168 508580 169174 508592
rect 508498 508580 508504 508592
rect 508556 508580 508562 508632
rect 7926 508512 7932 508564
rect 7984 508552 7990 508564
rect 354398 508552 354404 508564
rect 7984 508524 354404 508552
rect 7984 508512 7990 508524
rect 354398 508512 354404 508524
rect 354456 508512 354462 508564
rect 361114 508552 361120 508564
rect 354646 508524 361120 508552
rect 7834 508444 7840 508496
rect 7892 508484 7898 508496
rect 354646 508484 354674 508524
rect 361114 508512 361120 508524
rect 361172 508512 361178 508564
rect 356698 508484 356704 508496
rect 7892 508456 354674 508484
rect 356659 508456 356704 508484
rect 7892 508444 7898 508456
rect 356698 508444 356704 508456
rect 356756 508444 356762 508496
rect 358906 508484 358912 508496
rect 358867 508456 358912 508484
rect 358906 508444 358912 508456
rect 358964 508444 358970 508496
rect 363322 508484 363328 508496
rect 363283 508456 363328 508484
rect 363322 508444 363328 508456
rect 363380 508444 363386 508496
rect 220446 508376 220452 508428
rect 220504 508416 220510 508428
rect 573358 508416 573364 508428
rect 220504 508388 573364 508416
rect 220504 508376 220510 508388
rect 573358 508376 573364 508388
rect 573416 508376 573422 508428
rect 7742 508308 7748 508360
rect 7800 508348 7806 508360
rect 367830 508348 367836 508360
rect 7800 508320 367836 508348
rect 7800 508308 7806 508320
rect 367830 508308 367836 508320
rect 367888 508308 367894 508360
rect 370038 508348 370044 508360
rect 369999 508320 370044 508348
rect 370038 508308 370044 508320
rect 370096 508308 370102 508360
rect 9030 508240 9036 508292
rect 9088 508280 9094 508292
rect 374546 508280 374552 508292
rect 9088 508252 374552 508280
rect 9088 508240 9094 508252
rect 374546 508240 374552 508252
rect 374604 508240 374610 508292
rect 10502 508172 10508 508224
rect 10560 508212 10566 508224
rect 381262 508212 381268 508224
rect 10560 508184 381268 508212
rect 10560 508172 10566 508184
rect 381262 508172 381268 508184
rect 381320 508172 381326 508224
rect 383470 508212 383476 508224
rect 383431 508184 383476 508212
rect 383470 508172 383476 508184
rect 383528 508172 383534 508224
rect 8938 508104 8944 508156
rect 8996 508144 9002 508156
rect 387886 508144 387892 508156
rect 8996 508116 387892 508144
rect 8996 508104 9002 508116
rect 387886 508104 387892 508116
rect 387944 508104 387950 508156
rect 10410 508036 10416 508088
rect 10468 508076 10474 508088
rect 394602 508076 394608 508088
rect 10468 508048 394608 508076
rect 10468 508036 10474 508048
rect 394602 508036 394608 508048
rect 394660 508036 394666 508088
rect 401318 508076 401324 508088
rect 396368 508048 401324 508076
rect 7650 507968 7656 508020
rect 7708 508008 7714 508020
rect 396368 508008 396396 508048
rect 401318 508036 401324 508048
rect 401376 508036 401382 508088
rect 396534 508008 396540 508020
rect 7708 507980 396396 508008
rect 396495 507980 396540 508008
rect 7708 507968 7714 507980
rect 396534 507968 396540 507980
rect 396592 507968 396598 508020
rect 7558 507900 7564 507952
rect 7616 507940 7622 507952
rect 407758 507940 407764 507952
rect 7616 507912 407764 507940
rect 7616 507900 7622 507912
rect 407758 507900 407764 507912
rect 407816 507900 407822 507952
rect 10318 507832 10324 507884
rect 10376 507872 10382 507884
rect 414382 507872 414388 507884
rect 10376 507844 414388 507872
rect 10376 507832 10382 507844
rect 414382 507832 414388 507844
rect 414440 507832 414446 507884
rect 236362 507764 236368 507816
rect 236420 507804 236426 507816
rect 426066 507804 426072 507816
rect 236420 507776 426072 507804
rect 236420 507764 236426 507776
rect 426066 507764 426072 507776
rect 426124 507764 426130 507816
rect 211890 507696 211896 507748
rect 211948 507736 211954 507748
rect 211948 507708 219434 507736
rect 211948 507696 211954 507708
rect 218514 507668 218520 507680
rect 218475 507640 218520 507668
rect 218514 507628 218520 507640
rect 218572 507628 218578 507680
rect 219406 507668 219434 507708
rect 227530 507696 227536 507748
rect 227588 507736 227594 507748
rect 425974 507736 425980 507748
rect 227588 507708 425980 507736
rect 227588 507696 227594 507708
rect 425974 507696 425980 507708
rect 426032 507696 426038 507748
rect 429930 507668 429936 507680
rect 219406 507640 429936 507668
rect 429930 507628 429936 507640
rect 429988 507628 429994 507680
rect 205082 507600 205088 507612
rect 205043 507572 205088 507600
rect 205082 507560 205088 507572
rect 205140 507560 205146 507612
rect 209498 507560 209504 507612
rect 209556 507600 209562 507612
rect 430022 507600 430028 507612
rect 209556 507572 430028 507600
rect 209556 507560 209562 507572
rect 430022 507560 430028 507572
rect 430080 507560 430086 507612
rect 202782 507492 202788 507544
rect 202840 507532 202846 507544
rect 428734 507532 428740 507544
rect 202840 507504 428740 507532
rect 202840 507492 202846 507504
rect 428734 507492 428740 507504
rect 428792 507492 428798 507544
rect 195790 507424 195796 507476
rect 195848 507464 195854 507476
rect 428642 507464 428648 507476
rect 195848 507436 428648 507464
rect 195848 507424 195854 507436
rect 428642 507424 428648 507436
rect 428700 507424 428706 507476
rect 191650 507356 191656 507408
rect 191708 507396 191714 507408
rect 429838 507396 429844 507408
rect 191708 507368 429844 507396
rect 191708 507356 191714 507368
rect 429838 507356 429844 507368
rect 429896 507356 429902 507408
rect 182818 507288 182824 507340
rect 182876 507328 182882 507340
rect 182876 507300 186452 507328
rect 182876 507288 182882 507300
rect 184934 507220 184940 507272
rect 184992 507220 184998 507272
rect 186424 507260 186452 507300
rect 189442 507288 189448 507340
rect 189500 507328 189506 507340
rect 428550 507328 428556 507340
rect 189500 507300 428556 507328
rect 189500 507288 189506 507300
rect 428550 507288 428556 507300
rect 428608 507288 428614 507340
rect 349525 507263 349583 507269
rect 349525 507260 349537 507263
rect 186424 507232 349537 507260
rect 349525 507229 349537 507232
rect 349571 507229 349583 507263
rect 349525 507223 349583 507229
rect 349706 507220 349712 507272
rect 349764 507220 349770 507272
rect 349893 507263 349951 507269
rect 349893 507229 349905 507263
rect 349939 507260 349951 507263
rect 425790 507260 425796 507272
rect 349939 507232 425796 507260
rect 349939 507229 349951 507232
rect 349893 507223 349951 507229
rect 425790 507220 425796 507232
rect 425848 507220 425854 507272
rect 184952 507192 184980 507220
rect 349617 507195 349675 507201
rect 349617 507192 349629 507195
rect 184952 507164 349629 507192
rect 349617 507161 349629 507164
rect 349663 507161 349675 507195
rect 349617 507155 349675 507161
rect 237377 507127 237435 507133
rect 237377 507093 237389 507127
rect 237423 507124 237435 507127
rect 349525 507127 349583 507133
rect 349525 507124 349537 507127
rect 237423 507096 349537 507124
rect 237423 507093 237435 507096
rect 237377 507087 237435 507093
rect 349525 507093 349537 507096
rect 349571 507093 349583 507127
rect 349525 507087 349583 507093
rect 5534 507016 5540 507068
rect 5592 507056 5598 507068
rect 349724 507056 349752 507220
rect 349801 507195 349859 507201
rect 349801 507161 349813 507195
rect 349847 507192 349859 507195
rect 428458 507192 428464 507204
rect 349847 507164 428464 507192
rect 349847 507161 349859 507164
rect 349801 507155 349859 507161
rect 428458 507152 428464 507164
rect 428516 507152 428522 507204
rect 349893 507127 349951 507133
rect 349893 507093 349905 507127
rect 349939 507124 349951 507127
rect 580258 507124 580264 507136
rect 349939 507096 580264 507124
rect 349939 507093 349951 507096
rect 349893 507087 349951 507093
rect 580258 507084 580264 507096
rect 580316 507084 580322 507136
rect 5592 507028 349752 507056
rect 5592 507016 5598 507028
rect 11974 506948 11980 507000
rect 12032 506988 12038 507000
rect 356701 506991 356759 506997
rect 356701 506988 356713 506991
rect 12032 506960 356713 506988
rect 12032 506948 12038 506960
rect 356701 506957 356713 506960
rect 356747 506957 356759 506991
rect 356701 506951 356759 506957
rect 11882 506880 11888 506932
rect 11940 506920 11946 506932
rect 363325 506923 363383 506929
rect 363325 506920 363337 506923
rect 11940 506892 363337 506920
rect 11940 506880 11946 506892
rect 363325 506889 363337 506892
rect 363371 506889 363383 506923
rect 363325 506883 363383 506889
rect 5074 506812 5080 506864
rect 5132 506852 5138 506864
rect 358909 506855 358967 506861
rect 358909 506852 358921 506855
rect 5132 506824 358921 506852
rect 5132 506812 5138 506824
rect 358909 506821 358921 506824
rect 358955 506821 358967 506855
rect 358909 506815 358967 506821
rect 11790 506744 11796 506796
rect 11848 506784 11854 506796
rect 370041 506787 370099 506793
rect 370041 506784 370053 506787
rect 11848 506756 370053 506784
rect 11848 506744 11854 506756
rect 370041 506753 370053 506756
rect 370087 506753 370099 506787
rect 370041 506747 370099 506753
rect 218517 506719 218575 506725
rect 218517 506685 218529 506719
rect 218563 506716 218575 506719
rect 580442 506716 580448 506728
rect 218563 506688 580448 506716
rect 218563 506685 218575 506688
rect 218517 506679 218575 506685
rect 580442 506676 580448 506688
rect 580500 506676 580506 506728
rect 205085 506651 205143 506657
rect 205085 506617 205097 506651
rect 205131 506648 205143 506651
rect 580350 506648 580356 506660
rect 205131 506620 580356 506648
rect 205131 506617 205143 506620
rect 205085 506611 205143 506617
rect 580350 506608 580356 506620
rect 580408 506608 580414 506660
rect 3602 506540 3608 506592
rect 3660 506580 3666 506592
rect 383473 506583 383531 506589
rect 383473 506580 383485 506583
rect 3660 506552 383485 506580
rect 3660 506540 3666 506552
rect 383473 506549 383485 506552
rect 383519 506549 383531 506583
rect 383473 506543 383531 506549
rect 3510 506472 3516 506524
rect 3568 506512 3574 506524
rect 396537 506515 396595 506521
rect 396537 506512 396549 506515
rect 3568 506484 396549 506512
rect 3568 506472 3574 506484
rect 396537 506481 396549 506484
rect 396583 506481 396595 506515
rect 396537 506475 396595 506481
rect 3142 502256 3148 502308
rect 3200 502296 3206 502308
rect 5534 502296 5540 502308
rect 3200 502268 5540 502296
rect 3200 502256 3206 502268
rect 5534 502256 5540 502268
rect 5592 502256 5598 502308
rect 426066 485732 426072 485784
rect 426124 485772 426130 485784
rect 580166 485772 580172 485784
rect 426124 485744 580172 485772
rect 426124 485732 426130 485744
rect 580166 485732 580172 485744
rect 580224 485732 580230 485784
rect 3326 475668 3332 475720
rect 3384 475708 3390 475720
rect 7926 475708 7932 475720
rect 3384 475680 7932 475708
rect 3384 475668 3390 475680
rect 7926 475668 7932 475680
rect 7984 475668 7990 475720
rect 431310 471928 431316 471980
rect 431368 471968 431374 471980
rect 580166 471968 580172 471980
rect 431368 471940 580172 471968
rect 431368 471928 431374 471940
rect 580166 471928 580172 471940
rect 580224 471928 580230 471980
rect 2774 463428 2780 463480
rect 2832 463468 2838 463480
rect 5074 463468 5080 463480
rect 2832 463440 5080 463468
rect 2832 463428 2838 463440
rect 5074 463428 5080 463440
rect 5132 463428 5138 463480
rect 421926 458124 421932 458176
rect 421984 458164 421990 458176
rect 580166 458164 580172 458176
rect 421984 458136 580172 458164
rect 421984 458124 421990 458136
rect 580166 458124 580172 458136
rect 580224 458124 580230 458176
rect 3326 449828 3332 449880
rect 3384 449868 3390 449880
rect 11974 449868 11980 449880
rect 3384 449840 11980 449868
rect 3384 449828 3390 449840
rect 11974 449828 11980 449840
rect 12032 449828 12038 449880
rect 430114 431876 430120 431928
rect 430172 431916 430178 431928
rect 580166 431916 580172 431928
rect 430172 431888 580172 431916
rect 430172 431876 430178 431888
rect 580166 431876 580172 431888
rect 580224 431876 580230 431928
rect 3326 423580 3332 423632
rect 3384 423620 3390 423632
rect 7834 423620 7840 423632
rect 3384 423592 7840 423620
rect 3384 423580 3390 423592
rect 7834 423580 7840 423592
rect 7892 423580 7898 423632
rect 431218 419432 431224 419484
rect 431276 419472 431282 419484
rect 579706 419472 579712 419484
rect 431276 419444 579712 419472
rect 431276 419432 431282 419444
rect 579706 419432 579712 419444
rect 579764 419432 579770 419484
rect 2774 411000 2780 411052
rect 2832 411040 2838 411052
rect 4982 411040 4988 411052
rect 2832 411012 4988 411040
rect 2832 411000 2838 411012
rect 4982 411000 4988 411012
rect 5040 411000 5046 411052
rect 425974 405628 425980 405680
rect 426032 405668 426038 405680
rect 579798 405668 579804 405680
rect 426032 405640 579804 405668
rect 426032 405628 426038 405640
rect 579798 405628 579804 405640
rect 579856 405628 579862 405680
rect 3326 398760 3332 398812
rect 3384 398800 3390 398812
rect 11882 398800 11888 398812
rect 3384 398772 11888 398800
rect 3384 398760 3390 398772
rect 11882 398760 11888 398772
rect 11940 398760 11946 398812
rect 562318 379448 562324 379500
rect 562376 379488 562382 379500
rect 579798 379488 579804 379500
rect 562376 379460 579804 379488
rect 562376 379448 562382 379460
rect 579798 379448 579804 379460
rect 579856 379448 579862 379500
rect 3050 372376 3056 372428
rect 3108 372416 3114 372428
rect 7742 372416 7748 372428
rect 3108 372388 7748 372416
rect 3108 372376 3114 372388
rect 7742 372376 7748 372388
rect 7800 372376 7806 372428
rect 496078 365644 496084 365696
rect 496136 365684 496142 365696
rect 580166 365684 580172 365696
rect 496136 365656 580172 365684
rect 496136 365644 496142 365656
rect 580166 365644 580172 365656
rect 580224 365644 580230 365696
rect 2774 358436 2780 358488
rect 2832 358476 2838 358488
rect 4890 358476 4896 358488
rect 2832 358448 4896 358476
rect 2832 358436 2838 358448
rect 4890 358436 4896 358448
rect 4948 358436 4954 358488
rect 573358 353200 573364 353252
rect 573416 353240 573422 353252
rect 579614 353240 579620 353252
rect 573416 353212 579620 353240
rect 573416 353200 573422 353212
rect 579614 353200 579620 353212
rect 579672 353200 579678 353252
rect 3326 346332 3332 346384
rect 3384 346372 3390 346384
rect 11790 346372 11796 346384
rect 3384 346344 11796 346372
rect 3384 346332 3390 346344
rect 11790 346332 11796 346344
rect 11848 346332 11854 346384
rect 478138 325592 478144 325644
rect 478196 325632 478202 325644
rect 580166 325632 580172 325644
rect 478196 325604 580172 325632
rect 478196 325592 478202 325604
rect 580166 325592 580172 325604
rect 580224 325592 580230 325644
rect 3326 319540 3332 319592
rect 3384 319580 3390 319592
rect 9030 319580 9036 319592
rect 3384 319552 9036 319580
rect 3384 319540 3390 319552
rect 9030 319540 9036 319552
rect 9088 319540 9094 319592
rect 3326 306280 3332 306332
rect 3384 306320 3390 306332
rect 11698 306320 11704 306332
rect 3384 306292 11704 306320
rect 3384 306280 3390 306292
rect 11698 306280 11704 306292
rect 11756 306280 11762 306332
rect 425882 299412 425888 299464
rect 425940 299452 425946 299464
rect 580166 299452 580172 299464
rect 425940 299424 580172 299452
rect 425940 299412 425946 299424
rect 580166 299412 580172 299424
rect 580224 299412 580230 299464
rect 2866 293904 2872 293956
rect 2924 293944 2930 293956
rect 14642 293944 14648 293956
rect 2924 293916 14648 293944
rect 2924 293904 2930 293916
rect 14642 293904 14648 293916
rect 14700 293904 14706 293956
rect 430022 273164 430028 273216
rect 430080 273204 430086 273216
rect 580166 273204 580172 273216
rect 430080 273176 580172 273204
rect 430080 273164 430086 273176
rect 580166 273164 580172 273176
rect 580224 273164 580230 273216
rect 3234 267656 3240 267708
rect 3292 267696 3298 267708
rect 10502 267696 10508 267708
rect 3292 267668 10508 267696
rect 3292 267656 3298 267668
rect 10502 267656 10508 267668
rect 10560 267656 10566 267708
rect 429930 259360 429936 259412
rect 429988 259400 429994 259412
rect 579614 259400 579620 259412
rect 429988 259372 579620 259400
rect 429988 259360 429994 259372
rect 579614 259360 579620 259372
rect 579672 259360 579678 259412
rect 3326 255212 3332 255264
rect 3384 255252 3390 255264
rect 14550 255252 14556 255264
rect 3384 255224 14556 255252
rect 3384 255212 3390 255224
rect 14550 255212 14556 255224
rect 14608 255212 14614 255264
rect 424502 245556 424508 245608
rect 424560 245596 424566 245608
rect 580166 245596 580172 245608
rect 424560 245568 580172 245596
rect 424560 245556 424566 245568
rect 580166 245556 580172 245568
rect 580224 245556 580230 245608
rect 428734 233180 428740 233232
rect 428792 233220 428798 233232
rect 580166 233220 580172 233232
rect 428792 233192 580172 233220
rect 428792 233180 428798 233192
rect 580166 233180 580172 233192
rect 580224 233180 580230 233232
rect 3326 214956 3332 215008
rect 3384 214996 3390 215008
rect 8938 214996 8944 215008
rect 3384 214968 8944 214996
rect 3384 214956 3390 214968
rect 8938 214956 8944 214968
rect 8996 214956 9002 215008
rect 422938 206932 422944 206984
rect 422996 206972 423002 206984
rect 580166 206972 580172 206984
rect 422996 206944 580172 206972
rect 422996 206932 423002 206944
rect 580166 206932 580172 206944
rect 580224 206932 580230 206984
rect 3050 202784 3056 202836
rect 3108 202824 3114 202836
rect 14458 202824 14464 202836
rect 3108 202796 14464 202824
rect 3108 202784 3114 202796
rect 14458 202784 14464 202796
rect 14516 202784 14522 202836
rect 168466 200404 168472 200456
rect 168524 200444 168530 200456
rect 168742 200444 168748 200456
rect 168524 200416 168748 200444
rect 168524 200404 168530 200416
rect 168742 200404 168748 200416
rect 168800 200404 168806 200456
rect 240226 200404 240232 200456
rect 240284 200444 240290 200456
rect 240502 200444 240508 200456
rect 240284 200416 240508 200444
rect 240284 200404 240290 200416
rect 240502 200404 240508 200416
rect 240560 200404 240566 200456
rect 252554 200404 252560 200456
rect 252612 200444 252618 200456
rect 252830 200444 252836 200456
rect 252612 200416 252836 200444
rect 252612 200404 252618 200416
rect 252830 200404 252836 200416
rect 252888 200404 252894 200456
rect 61378 198636 61384 198688
rect 61436 198676 61442 198688
rect 174446 198676 174452 198688
rect 61436 198648 174452 198676
rect 61436 198636 61442 198648
rect 174446 198636 174452 198648
rect 174504 198636 174510 198688
rect 177298 198636 177304 198688
rect 177356 198676 177362 198688
rect 218146 198676 218152 198688
rect 177356 198648 218152 198676
rect 177356 198636 177362 198648
rect 218146 198636 218152 198648
rect 218204 198636 218210 198688
rect 238662 198636 238668 198688
rect 238720 198676 238726 198688
rect 269390 198676 269396 198688
rect 238720 198648 269396 198676
rect 238720 198636 238726 198648
rect 269390 198636 269396 198648
rect 269448 198636 269454 198688
rect 277302 198636 277308 198688
rect 277360 198676 277366 198688
rect 285950 198676 285956 198688
rect 277360 198648 285956 198676
rect 277360 198636 277366 198648
rect 285950 198636 285956 198648
rect 286008 198636 286014 198688
rect 312906 198636 312912 198688
rect 312964 198676 312970 198688
rect 335538 198676 335544 198688
rect 312964 198648 335544 198676
rect 312964 198636 312970 198648
rect 335538 198636 335544 198648
rect 335596 198636 335602 198688
rect 337930 198636 337936 198688
rect 337988 198676 337994 198688
rect 393498 198676 393504 198688
rect 337988 198648 393504 198676
rect 337988 198636 337994 198648
rect 393498 198636 393504 198648
rect 393556 198636 393562 198688
rect 395522 198636 395528 198688
rect 395580 198676 395586 198688
rect 400033 198679 400091 198685
rect 400033 198676 400045 198679
rect 395580 198648 400045 198676
rect 395580 198636 395586 198648
rect 400033 198645 400045 198648
rect 400079 198645 400091 198679
rect 400033 198639 400091 198645
rect 400122 198636 400128 198688
rect 400180 198676 400186 198688
rect 471238 198676 471244 198688
rect 400180 198648 471244 198676
rect 400180 198636 400186 198648
rect 471238 198636 471244 198648
rect 471296 198636 471302 198688
rect 76558 198568 76564 198620
rect 76616 198608 76622 198620
rect 195054 198608 195060 198620
rect 76616 198580 195060 198608
rect 76616 198568 76622 198580
rect 195054 198568 195060 198580
rect 195112 198568 195118 198620
rect 196894 198568 196900 198620
rect 196952 198608 196958 198620
rect 213086 198608 213092 198620
rect 196952 198580 213092 198608
rect 196952 198568 196958 198580
rect 213086 198568 213092 198580
rect 213144 198568 213150 198620
rect 213270 198568 213276 198620
rect 213328 198608 213334 198620
rect 229646 198608 229652 198620
rect 213328 198580 229652 198608
rect 213328 198568 213334 198580
rect 229646 198568 229652 198580
rect 229704 198568 229710 198620
rect 235902 198568 235908 198620
rect 235960 198608 235966 198620
rect 267918 198608 267924 198620
rect 235960 198580 267924 198608
rect 235960 198568 235966 198580
rect 267918 198568 267924 198580
rect 267976 198568 267982 198620
rect 271782 198568 271788 198620
rect 271840 198608 271846 198620
rect 283926 198608 283932 198620
rect 271840 198580 283932 198608
rect 271840 198568 271846 198580
rect 283926 198568 283932 198580
rect 283984 198568 283990 198620
rect 319162 198568 319168 198620
rect 319220 198608 319226 198620
rect 335998 198608 336004 198620
rect 319220 198580 336004 198608
rect 319220 198568 319226 198580
rect 335998 198568 336004 198580
rect 336056 198568 336062 198620
rect 347498 198568 347504 198620
rect 347556 198608 347562 198620
rect 414566 198608 414572 198620
rect 347556 198580 414572 198608
rect 347556 198568 347562 198580
rect 414566 198568 414572 198580
rect 414624 198568 414630 198620
rect 419350 198568 419356 198620
rect 419408 198608 419414 198620
rect 490558 198608 490564 198620
rect 419408 198580 490564 198608
rect 419408 198568 419414 198580
rect 490558 198568 490564 198580
rect 490616 198568 490622 198620
rect 71038 198500 71044 198552
rect 71096 198540 71102 198552
rect 191926 198540 191932 198552
rect 71096 198512 191932 198540
rect 71096 198500 71102 198512
rect 191926 198500 191932 198512
rect 191984 198500 191990 198552
rect 197998 198500 198004 198552
rect 198056 198540 198062 198552
rect 214742 198540 214748 198552
rect 198056 198512 214748 198540
rect 198056 198500 198062 198512
rect 214742 198500 214748 198512
rect 214800 198500 214806 198552
rect 217318 198500 217324 198552
rect 217376 198540 217382 198552
rect 227714 198540 227720 198552
rect 217376 198512 227720 198540
rect 217376 198500 217382 198512
rect 227714 198500 227720 198512
rect 227772 198500 227778 198552
rect 234522 198500 234528 198552
rect 234580 198540 234586 198552
rect 267366 198540 267372 198552
rect 234580 198512 267372 198540
rect 234580 198500 234586 198512
rect 267366 198500 267372 198512
rect 267424 198500 267430 198552
rect 269022 198500 269028 198552
rect 269080 198540 269086 198552
rect 282270 198540 282276 198552
rect 269080 198512 282276 198540
rect 269080 198500 269086 198512
rect 282270 198500 282276 198512
rect 282328 198500 282334 198552
rect 298370 198500 298376 198552
rect 298428 198540 298434 198552
rect 302510 198540 302516 198552
rect 298428 198512 302516 198540
rect 298428 198500 298434 198512
rect 302510 198500 302516 198512
rect 302568 198500 302574 198552
rect 311802 198500 311808 198552
rect 311860 198540 311866 198552
rect 330478 198540 330484 198552
rect 311860 198512 330484 198540
rect 311860 198500 311866 198512
rect 330478 198500 330484 198512
rect 330536 198500 330542 198552
rect 332962 198500 332968 198552
rect 333020 198540 333026 198552
rect 340230 198540 340236 198552
rect 333020 198512 340236 198540
rect 333020 198500 333026 198512
rect 340230 198500 340236 198512
rect 340288 198500 340294 198552
rect 350442 198500 350448 198552
rect 350500 198540 350506 198552
rect 420181 198543 420239 198549
rect 420181 198540 420193 198543
rect 350500 198512 420193 198540
rect 350500 198500 350506 198512
rect 420181 198509 420193 198512
rect 420227 198509 420239 198543
rect 420181 198503 420239 198509
rect 420362 198500 420368 198552
rect 420420 198540 420426 198552
rect 420822 198540 420828 198552
rect 420420 198512 420828 198540
rect 420420 198500 420426 198512
rect 420822 198500 420828 198512
rect 420880 198500 420886 198552
rect 58618 198432 58624 198484
rect 58676 198472 58682 198484
rect 184198 198472 184204 198484
rect 58676 198444 184204 198472
rect 58676 198432 58682 198444
rect 184198 198432 184204 198444
rect 184256 198432 184262 198484
rect 184290 198432 184296 198484
rect 184348 198472 184354 198484
rect 193582 198472 193588 198484
rect 184348 198444 193588 198472
rect 184348 198432 184354 198444
rect 193582 198432 193588 198444
rect 193640 198432 193646 198484
rect 195238 198432 195244 198484
rect 195296 198472 195302 198484
rect 201681 198475 201739 198481
rect 195296 198444 201632 198472
rect 195296 198432 195302 198444
rect 51718 198364 51724 198416
rect 51776 198404 51782 198416
rect 181070 198404 181076 198416
rect 51776 198376 181076 198404
rect 51776 198364 51782 198376
rect 181070 198364 181076 198376
rect 181128 198364 181134 198416
rect 185578 198364 185584 198416
rect 185636 198404 185642 198416
rect 196526 198404 196532 198416
rect 185636 198376 196532 198404
rect 185636 198364 185642 198376
rect 196526 198364 196532 198376
rect 196584 198364 196590 198416
rect 201497 198407 201555 198413
rect 201497 198404 201509 198407
rect 196636 198376 201509 198404
rect 57238 198296 57244 198348
rect 57296 198336 57302 198348
rect 189074 198336 189080 198348
rect 57296 198308 189080 198336
rect 57296 198296 57302 198308
rect 189074 198296 189080 198308
rect 189132 198296 189138 198348
rect 193858 198296 193864 198348
rect 193916 198336 193922 198348
rect 196636 198336 196664 198376
rect 201497 198373 201509 198376
rect 201543 198373 201555 198407
rect 201604 198404 201632 198444
rect 201681 198441 201693 198475
rect 201727 198472 201739 198475
rect 214006 198472 214012 198484
rect 201727 198444 214012 198472
rect 201727 198441 201739 198444
rect 201681 198435 201739 198441
rect 214006 198432 214012 198444
rect 214064 198432 214070 198484
rect 214650 198432 214656 198484
rect 214708 198472 214714 198484
rect 226518 198472 226524 198484
rect 214708 198444 226524 198472
rect 214708 198432 214714 198444
rect 226518 198432 226524 198444
rect 226576 198432 226582 198484
rect 231762 198432 231768 198484
rect 231820 198472 231826 198484
rect 266354 198472 266360 198484
rect 231820 198444 266360 198472
rect 231820 198432 231826 198444
rect 266354 198432 266360 198444
rect 266412 198432 266418 198484
rect 270402 198432 270408 198484
rect 270460 198472 270466 198484
rect 283374 198472 283380 198484
rect 270460 198444 283380 198472
rect 270460 198432 270466 198444
rect 283374 198432 283380 198444
rect 283432 198432 283438 198484
rect 320082 198432 320088 198484
rect 320140 198472 320146 198484
rect 338758 198472 338764 198484
rect 320140 198444 338764 198472
rect 320140 198432 320146 198444
rect 338758 198432 338764 198444
rect 338816 198432 338822 198484
rect 353754 198432 353760 198484
rect 353812 198472 353818 198484
rect 429194 198472 429200 198484
rect 353812 198444 429200 198472
rect 353812 198432 353818 198444
rect 429194 198432 429200 198444
rect 429252 198432 429258 198484
rect 216766 198404 216772 198416
rect 201604 198376 216772 198404
rect 201497 198367 201555 198373
rect 216766 198364 216772 198376
rect 216824 198364 216830 198416
rect 227622 198364 227628 198416
rect 227680 198404 227686 198416
rect 264974 198404 264980 198416
rect 227680 198376 264980 198404
rect 227680 198364 227686 198376
rect 264974 198364 264980 198376
rect 265032 198364 265038 198416
rect 267642 198364 267648 198416
rect 267700 198404 267706 198416
rect 281718 198404 281724 198416
rect 267700 198376 281724 198404
rect 267700 198364 267706 198376
rect 281718 198364 281724 198376
rect 281776 198364 281782 198416
rect 299290 198364 299296 198416
rect 299348 198404 299354 198416
rect 305178 198404 305184 198416
rect 299348 198376 305184 198404
rect 299348 198364 299354 198376
rect 305178 198364 305184 198376
rect 305236 198364 305242 198416
rect 344370 198364 344376 198416
rect 344428 198404 344434 198416
rect 352558 198404 352564 198416
rect 344428 198376 352564 198404
rect 344428 198364 344434 198376
rect 352558 198364 352564 198376
rect 352616 198364 352622 198416
rect 356882 198364 356888 198416
rect 356940 198404 356946 198416
rect 436094 198404 436100 198416
rect 356940 198376 436100 198404
rect 356940 198364 356946 198376
rect 436094 198364 436100 198376
rect 436152 198364 436158 198416
rect 193916 198308 196664 198336
rect 193916 198296 193922 198308
rect 196802 198296 196808 198348
rect 196860 198336 196866 198348
rect 218238 198336 218244 198348
rect 196860 198308 218244 198336
rect 196860 198296 196866 198308
rect 218238 198296 218244 198308
rect 218296 198296 218302 198348
rect 223482 198296 223488 198348
rect 223540 198336 223546 198348
rect 262766 198336 262772 198348
rect 223540 198308 262772 198336
rect 223540 198296 223546 198308
rect 262766 198296 262772 198308
rect 262824 198296 262830 198348
rect 268930 198296 268936 198348
rect 268988 198336 268994 198348
rect 282914 198336 282920 198348
rect 268988 198308 282920 198336
rect 268988 198296 268994 198308
rect 282914 198296 282920 198308
rect 282972 198296 282978 198348
rect 326890 198296 326896 198348
rect 326948 198336 326954 198348
rect 353938 198336 353944 198348
rect 326948 198308 353944 198336
rect 326948 198296 326954 198308
rect 353938 198296 353944 198308
rect 353996 198296 354002 198348
rect 354646 198308 358308 198336
rect 35158 198228 35164 198280
rect 35216 198268 35222 198280
rect 178034 198268 178040 198280
rect 35216 198240 178040 198268
rect 35216 198228 35222 198240
rect 178034 198228 178040 198240
rect 178092 198228 178098 198280
rect 178678 198228 178684 198280
rect 178736 198268 178742 198280
rect 219434 198268 219440 198280
rect 178736 198240 219440 198268
rect 178736 198228 178742 198240
rect 219434 198228 219440 198240
rect 219492 198228 219498 198280
rect 220722 198228 220728 198280
rect 220780 198268 220786 198280
rect 261662 198268 261668 198280
rect 220780 198240 261668 198268
rect 220780 198228 220786 198240
rect 261662 198228 261668 198240
rect 261720 198228 261726 198280
rect 264882 198228 264888 198280
rect 264940 198268 264946 198280
rect 280798 198268 280804 198280
rect 264940 198240 280804 198268
rect 264940 198228 264946 198240
rect 280798 198228 280804 198240
rect 280856 198228 280862 198280
rect 285582 198228 285588 198280
rect 285640 198268 285646 198280
rect 290090 198268 290096 198280
rect 285640 198240 290096 198268
rect 285640 198228 285646 198240
rect 290090 198228 290096 198240
rect 290148 198228 290154 198280
rect 315942 198228 315948 198280
rect 316000 198268 316006 198280
rect 327902 198268 327908 198280
rect 316000 198240 327908 198268
rect 316000 198228 316006 198240
rect 327902 198228 327908 198240
rect 327960 198228 327966 198280
rect 330938 198228 330944 198280
rect 330996 198268 331002 198280
rect 354646 198268 354674 198308
rect 330996 198240 354674 198268
rect 330996 198228 331002 198240
rect 355778 198228 355784 198280
rect 355836 198268 355842 198280
rect 358170 198268 358176 198280
rect 355836 198240 358176 198268
rect 355836 198228 355842 198240
rect 358170 198228 358176 198240
rect 358228 198228 358234 198280
rect 358280 198268 358308 198308
rect 359826 198296 359832 198348
rect 359884 198336 359890 198348
rect 442994 198336 443000 198348
rect 359884 198308 443000 198336
rect 359884 198296 359890 198308
rect 442994 198296 443000 198308
rect 443052 198296 443058 198348
rect 361022 198268 361028 198280
rect 358280 198240 361028 198268
rect 361022 198228 361028 198240
rect 361080 198228 361086 198280
rect 362862 198228 362868 198280
rect 362920 198268 362926 198280
rect 449894 198268 449900 198280
rect 362920 198240 449900 198268
rect 362920 198228 362926 198240
rect 449894 198228 449900 198240
rect 449952 198228 449958 198280
rect 29638 198160 29644 198212
rect 29696 198200 29702 198212
rect 173986 198200 173992 198212
rect 29696 198172 173992 198200
rect 29696 198160 29702 198172
rect 173986 198160 173992 198172
rect 174044 198160 174050 198212
rect 184382 198160 184388 198212
rect 184440 198200 184446 198212
rect 216214 198200 216220 198212
rect 184440 198172 216220 198200
rect 184440 198160 184446 198172
rect 216214 198160 216220 198172
rect 216272 198160 216278 198212
rect 217962 198160 217968 198212
rect 218020 198200 218026 198212
rect 260190 198200 260196 198212
rect 218020 198172 260196 198200
rect 218020 198160 218026 198172
rect 260190 198160 260196 198172
rect 260248 198160 260254 198212
rect 262950 198160 262956 198212
rect 263008 198200 263014 198212
rect 279694 198200 279700 198212
rect 263008 198172 279700 198200
rect 263008 198160 263014 198172
rect 279694 198160 279700 198172
rect 279752 198160 279758 198212
rect 304074 198160 304080 198212
rect 304132 198200 304138 198212
rect 312538 198200 312544 198212
rect 304132 198172 312544 198200
rect 304132 198160 304138 198172
rect 312538 198160 312544 198172
rect 312596 198160 312602 198212
rect 318518 198160 318524 198212
rect 318576 198200 318582 198212
rect 349338 198200 349344 198212
rect 318576 198172 349344 198200
rect 318576 198160 318582 198172
rect 349338 198160 349344 198172
rect 349396 198160 349402 198212
rect 351822 198160 351828 198212
rect 351880 198200 351886 198212
rect 359458 198200 359464 198212
rect 351880 198172 359464 198200
rect 351880 198160 351886 198172
rect 359458 198160 359464 198172
rect 359516 198160 359522 198212
rect 359568 198172 364334 198200
rect 18598 198092 18604 198144
rect 18656 198132 18662 198144
rect 170214 198132 170220 198144
rect 18656 198104 170220 198132
rect 18656 198092 18662 198104
rect 170214 198092 170220 198104
rect 170272 198092 170278 198144
rect 191098 198092 191104 198144
rect 191156 198132 191162 198144
rect 207382 198132 207388 198144
rect 191156 198104 207388 198132
rect 191156 198092 191162 198104
rect 207382 198092 207388 198104
rect 207440 198092 207446 198144
rect 213822 198092 213828 198144
rect 213880 198132 213886 198144
rect 258534 198132 258540 198144
rect 213880 198104 258540 198132
rect 213880 198092 213886 198104
rect 258534 198092 258540 198104
rect 258592 198092 258598 198144
rect 260650 198092 260656 198144
rect 260708 198132 260714 198144
rect 278774 198132 278780 198144
rect 260708 198104 278780 198132
rect 260708 198092 260714 198104
rect 278774 198092 278780 198104
rect 278832 198092 278838 198144
rect 285490 198092 285496 198144
rect 285548 198132 285554 198144
rect 289814 198132 289820 198144
rect 285548 198104 289820 198132
rect 285548 198092 285554 198104
rect 289814 198092 289820 198104
rect 289872 198092 289878 198144
rect 309778 198092 309784 198144
rect 309836 198132 309842 198144
rect 310422 198132 310428 198144
rect 309836 198104 310428 198132
rect 309836 198092 309842 198104
rect 310422 198092 310428 198104
rect 310480 198092 310486 198144
rect 323118 198132 323124 198144
rect 316006 198104 323124 198132
rect 11698 198024 11704 198076
rect 11756 198064 11762 198076
rect 167638 198064 167644 198076
rect 11756 198036 167644 198064
rect 11756 198024 11762 198036
rect 167638 198024 167644 198036
rect 167696 198024 167702 198076
rect 184198 198024 184204 198076
rect 184256 198064 184262 198076
rect 190454 198064 190460 198076
rect 184256 198036 190460 198064
rect 184256 198024 184262 198036
rect 190454 198024 190460 198036
rect 190512 198024 190518 198076
rect 192478 198024 192484 198076
rect 192536 198064 192542 198076
rect 210510 198064 210516 198076
rect 192536 198036 210516 198064
rect 192536 198024 192542 198036
rect 210510 198024 210516 198036
rect 210568 198024 210574 198076
rect 210970 198024 210976 198076
rect 211028 198064 211034 198076
rect 257062 198064 257068 198076
rect 211028 198036 257068 198064
rect 211028 198024 211034 198036
rect 257062 198024 257068 198036
rect 257120 198024 257126 198076
rect 259362 198024 259368 198076
rect 259420 198064 259426 198076
rect 278222 198064 278228 198076
rect 259420 198036 278228 198064
rect 259420 198024 259426 198036
rect 278222 198024 278228 198036
rect 278280 198024 278286 198076
rect 278682 198024 278688 198076
rect 278740 198064 278746 198076
rect 287054 198064 287060 198076
rect 278740 198036 287060 198064
rect 278740 198024 278746 198036
rect 287054 198024 287060 198036
rect 287112 198024 287118 198076
rect 302602 198024 302608 198076
rect 302660 198064 302666 198076
rect 311986 198064 311992 198076
rect 302660 198036 311992 198064
rect 302660 198024 302666 198036
rect 311986 198024 311992 198036
rect 312044 198024 312050 198076
rect 316006 198064 316034 198104
rect 323118 198092 323124 198104
rect 323176 198092 323182 198144
rect 327442 198092 327448 198144
rect 327500 198132 327506 198144
rect 358814 198132 358820 198144
rect 327500 198104 358820 198132
rect 327500 198092 327506 198104
rect 358814 198092 358820 198104
rect 358872 198092 358878 198144
rect 312096 198036 316034 198064
rect 14458 197956 14464 198008
rect 14516 197996 14522 198008
rect 169754 197996 169760 198008
rect 14516 197968 169760 197996
rect 14516 197956 14522 197968
rect 169754 197956 169760 197968
rect 169812 197956 169818 198008
rect 170398 197956 170404 198008
rect 170456 197996 170462 198008
rect 180794 197996 180800 198008
rect 170456 197968 180800 197996
rect 170456 197956 170462 197968
rect 180794 197956 180800 197968
rect 180852 197956 180858 198008
rect 182818 197956 182824 198008
rect 182876 197996 182882 198008
rect 187326 197996 187332 198008
rect 182876 197968 187332 197996
rect 182876 197956 182882 197968
rect 187326 197956 187332 197968
rect 187384 197956 187390 198008
rect 189718 197956 189724 198008
rect 189776 197996 189782 198008
rect 204254 197996 204260 198008
rect 189776 197968 204260 197996
rect 189776 197956 189782 197968
rect 204254 197956 204260 197968
rect 204312 197956 204318 198008
rect 206922 197956 206928 198008
rect 206980 197996 206986 198008
rect 255406 197996 255412 198008
rect 206980 197968 255412 197996
rect 206980 197956 206986 197968
rect 255406 197956 255412 197968
rect 255464 197956 255470 198008
rect 255958 197956 255964 198008
rect 256016 197996 256022 198008
rect 275646 197996 275652 198008
rect 256016 197968 275652 197996
rect 256016 197956 256022 197968
rect 275646 197956 275652 197968
rect 275704 197956 275710 198008
rect 276658 197956 276664 198008
rect 276716 197996 276722 198008
rect 285674 197996 285680 198008
rect 276716 197968 285680 197996
rect 276716 197956 276722 197968
rect 285674 197956 285680 197968
rect 285732 197956 285738 198008
rect 286962 197956 286968 198008
rect 287020 197996 287026 198008
rect 290550 197996 290556 198008
rect 287020 197968 290556 197996
rect 287020 197956 287026 197968
rect 290550 197956 290556 197968
rect 290608 197956 290614 198008
rect 295794 197956 295800 198008
rect 295852 197996 295858 198008
rect 296622 197996 296628 198008
rect 295852 197968 296628 197996
rect 295852 197956 295858 197968
rect 296622 197956 296628 197968
rect 296680 197956 296686 198008
rect 307202 197956 307208 198008
rect 307260 197996 307266 198008
rect 312096 197996 312124 198036
rect 317322 198024 317328 198076
rect 317380 198064 317386 198076
rect 318058 198064 318064 198076
rect 317380 198036 318064 198064
rect 317380 198024 317386 198036
rect 318058 198024 318064 198036
rect 318116 198024 318122 198076
rect 357802 198024 357808 198076
rect 357860 198064 357866 198076
rect 359568 198064 359596 198172
rect 363690 198132 363696 198144
rect 357860 198036 359596 198064
rect 359660 198104 363696 198132
rect 357860 198024 357866 198036
rect 307260 197968 312124 197996
rect 307260 197956 307266 197968
rect 314010 197956 314016 198008
rect 314068 197996 314074 198008
rect 314562 197996 314568 198008
rect 314068 197968 314568 197996
rect 314068 197956 314074 197968
rect 314562 197956 314568 197968
rect 314620 197956 314626 198008
rect 327718 197996 327724 198008
rect 316006 197968 327724 197996
rect 94498 197888 94504 197940
rect 94556 197928 94562 197940
rect 205910 197928 205916 197940
rect 94556 197900 205916 197928
rect 94556 197888 94562 197900
rect 205910 197888 205916 197900
rect 205968 197888 205974 197940
rect 209038 197888 209044 197940
rect 209096 197928 209102 197940
rect 241054 197928 241060 197940
rect 209096 197900 241060 197928
rect 209096 197888 209102 197900
rect 241054 197888 241060 197900
rect 241112 197888 241118 197940
rect 241422 197888 241428 197940
rect 241480 197928 241486 197940
rect 270586 197928 270592 197940
rect 241480 197900 270592 197928
rect 241480 197888 241486 197900
rect 270586 197888 270592 197900
rect 270644 197888 270650 197940
rect 310330 197888 310336 197940
rect 310388 197928 310394 197940
rect 316006 197928 316034 197968
rect 327718 197956 327724 197968
rect 327776 197956 327782 198008
rect 329742 197956 329748 198008
rect 329800 197996 329806 198008
rect 359660 197996 359688 198104
rect 363690 198092 363696 198104
rect 363748 198092 363754 198144
rect 364306 198132 364334 198172
rect 366910 198160 366916 198212
rect 366968 198200 366974 198212
rect 385586 198200 385592 198212
rect 366968 198172 385592 198200
rect 366968 198160 366974 198172
rect 385586 198160 385592 198172
rect 385644 198160 385650 198212
rect 392394 198160 392400 198212
rect 392452 198200 392458 198212
rect 482370 198200 482376 198212
rect 392452 198172 482376 198200
rect 392452 198160 392458 198172
rect 482370 198160 482376 198172
rect 482428 198160 482434 198212
rect 370590 198132 370596 198144
rect 364306 198104 370596 198132
rect 370590 198092 370596 198104
rect 370648 198092 370654 198144
rect 456794 198132 456800 198144
rect 370700 198104 456800 198132
rect 366082 198024 366088 198076
rect 366140 198064 366146 198076
rect 370700 198064 370728 198104
rect 456794 198092 456800 198104
rect 456852 198092 456858 198144
rect 366140 198036 370728 198064
rect 366140 198024 366146 198036
rect 370866 198024 370872 198076
rect 370924 198064 370930 198076
rect 467834 198064 467840 198076
rect 370924 198036 467840 198064
rect 370924 198024 370930 198036
rect 467834 198024 467840 198036
rect 467892 198024 467898 198076
rect 329800 197968 359688 197996
rect 329800 197956 329806 197968
rect 360930 197956 360936 198008
rect 360988 197996 360994 198008
rect 371970 197996 371976 198008
rect 360988 197968 371976 197996
rect 360988 197956 360994 197968
rect 371970 197956 371976 197968
rect 372028 197956 372034 198008
rect 373810 197956 373816 198008
rect 373868 197996 373874 198008
rect 474734 197996 474740 198008
rect 373868 197968 474740 197996
rect 373868 197956 373874 197968
rect 474734 197956 474740 197968
rect 474792 197956 474798 198008
rect 310388 197900 316034 197928
rect 310388 197888 310394 197900
rect 339218 197888 339224 197940
rect 339276 197928 339282 197940
rect 367738 197928 367744 197940
rect 339276 197900 367744 197928
rect 339276 197888 339282 197900
rect 367738 197888 367744 197900
rect 367796 197888 367802 197940
rect 369210 197888 369216 197940
rect 369268 197928 369274 197940
rect 393958 197928 393964 197940
rect 369268 197900 393964 197928
rect 369268 197888 369274 197900
rect 393958 197888 393964 197900
rect 394016 197888 394022 197940
rect 403618 197928 403624 197940
rect 396000 197900 403624 197928
rect 101582 197820 101588 197872
rect 101640 197860 101646 197872
rect 208946 197860 208952 197872
rect 101640 197832 208952 197860
rect 101640 197820 101646 197832
rect 208946 197820 208952 197832
rect 209004 197820 209010 197872
rect 209130 197820 209136 197872
rect 209188 197860 209194 197872
rect 239398 197860 239404 197872
rect 209188 197832 239404 197860
rect 209188 197820 209194 197832
rect 239398 197820 239404 197832
rect 239456 197820 239462 197872
rect 253842 197820 253848 197872
rect 253900 197860 253906 197872
rect 276198 197860 276204 197872
rect 253900 197832 276204 197860
rect 253900 197820 253906 197832
rect 276198 197820 276204 197832
rect 276256 197820 276262 197872
rect 298002 197820 298008 197872
rect 298060 197860 298066 197872
rect 298738 197860 298744 197872
rect 298060 197832 298744 197860
rect 298060 197820 298066 197832
rect 298738 197820 298744 197832
rect 298796 197820 298802 197872
rect 322106 197820 322112 197872
rect 322164 197860 322170 197872
rect 322842 197860 322848 197872
rect 322164 197832 322848 197860
rect 322164 197820 322170 197832
rect 322842 197820 322848 197832
rect 322900 197820 322906 197872
rect 328914 197820 328920 197872
rect 328972 197860 328978 197872
rect 329742 197860 329748 197872
rect 328972 197832 329748 197860
rect 328972 197820 328978 197832
rect 329742 197820 329748 197832
rect 329800 197820 329806 197872
rect 333514 197820 333520 197872
rect 333572 197860 333578 197872
rect 360930 197860 360936 197872
rect 333572 197832 360936 197860
rect 333572 197820 333578 197832
rect 360930 197820 360936 197832
rect 360988 197820 360994 197872
rect 367554 197820 367560 197872
rect 367612 197860 367618 197872
rect 367612 197832 367968 197860
rect 367612 197820 367618 197832
rect 107562 197752 107568 197804
rect 107620 197792 107626 197804
rect 212166 197792 212172 197804
rect 107620 197764 212172 197792
rect 107620 197752 107626 197764
rect 212166 197752 212172 197764
rect 212224 197752 212230 197804
rect 214558 197752 214564 197804
rect 214616 197792 214622 197804
rect 225046 197792 225052 197804
rect 214616 197764 225052 197792
rect 214616 197752 214622 197764
rect 225046 197752 225052 197764
rect 225104 197752 225110 197804
rect 232498 197752 232504 197804
rect 232556 197792 232562 197804
rect 261110 197792 261116 197804
rect 232556 197764 261116 197792
rect 232556 197752 232562 197764
rect 261110 197752 261116 197764
rect 261168 197752 261174 197804
rect 268378 197752 268384 197804
rect 268436 197792 268442 197804
rect 277670 197792 277676 197804
rect 268436 197764 277676 197792
rect 268436 197752 268442 197764
rect 277670 197752 277676 197764
rect 277728 197752 277734 197804
rect 326338 197752 326344 197804
rect 326396 197792 326402 197804
rect 340138 197792 340144 197804
rect 326396 197764 340144 197792
rect 326396 197752 326402 197764
rect 340138 197752 340144 197764
rect 340196 197752 340202 197804
rect 342162 197752 342168 197804
rect 342220 197792 342226 197804
rect 367830 197792 367836 197804
rect 342220 197764 367836 197792
rect 342220 197752 342226 197764
rect 367830 197752 367836 197764
rect 367888 197752 367894 197804
rect 367940 197792 367968 197832
rect 370130 197820 370136 197872
rect 370188 197860 370194 197872
rect 394881 197863 394939 197869
rect 394881 197860 394893 197863
rect 370188 197832 394893 197860
rect 370188 197820 370194 197832
rect 394881 197829 394893 197832
rect 394927 197829 394939 197863
rect 394881 197823 394939 197829
rect 394970 197820 394976 197872
rect 395028 197860 395034 197872
rect 395890 197860 395896 197872
rect 395028 197832 395896 197860
rect 395028 197820 395034 197832
rect 395890 197820 395896 197832
rect 395948 197820 395954 197872
rect 378778 197792 378784 197804
rect 367940 197764 378784 197792
rect 378778 197752 378784 197764
rect 378836 197752 378842 197804
rect 396000 197792 396028 197900
rect 403618 197888 403624 197900
rect 403676 197888 403682 197940
rect 407761 197931 407819 197937
rect 407761 197897 407773 197931
rect 407807 197928 407819 197931
rect 467098 197928 467104 197940
rect 407807 197900 467104 197928
rect 407807 197897 407819 197900
rect 407761 197891 407819 197897
rect 467098 197888 467104 197900
rect 467156 197888 467162 197940
rect 396994 197820 397000 197872
rect 397052 197860 397058 197872
rect 397052 197832 402974 197860
rect 397052 197820 397058 197832
rect 378888 197764 396028 197792
rect 397089 197795 397147 197801
rect 114462 197684 114468 197736
rect 114520 197724 114526 197736
rect 215294 197724 215300 197736
rect 114520 197696 215300 197724
rect 114520 197684 114526 197696
rect 215294 197684 215300 197696
rect 215352 197684 215358 197736
rect 216030 197684 216036 197736
rect 216088 197724 216094 197736
rect 236270 197724 236276 197736
rect 216088 197696 236276 197724
rect 216088 197684 216094 197696
rect 236270 197684 236276 197696
rect 236328 197684 236334 197736
rect 251818 197684 251824 197736
rect 251876 197724 251882 197736
rect 272518 197724 272524 197736
rect 251876 197696 272524 197724
rect 251876 197684 251882 197696
rect 272518 197684 272524 197696
rect 272576 197684 272582 197736
rect 306650 197684 306656 197736
rect 306708 197724 306714 197736
rect 307662 197724 307668 197736
rect 306708 197696 307668 197724
rect 306708 197684 306714 197696
rect 307662 197684 307668 197696
rect 307720 197684 307726 197736
rect 310882 197684 310888 197736
rect 310940 197724 310946 197736
rect 311802 197724 311808 197736
rect 310940 197696 311808 197724
rect 310940 197684 310946 197696
rect 311802 197684 311808 197696
rect 311860 197684 311866 197736
rect 320634 197684 320640 197736
rect 320692 197724 320698 197736
rect 321462 197724 321468 197736
rect 320692 197696 321468 197724
rect 320692 197684 320698 197696
rect 321462 197684 321468 197696
rect 321520 197684 321526 197736
rect 328270 197684 328276 197736
rect 328328 197724 328334 197736
rect 341518 197724 341524 197736
rect 328328 197696 341524 197724
rect 328328 197684 328334 197696
rect 341518 197684 341524 197696
rect 341576 197684 341582 197736
rect 343266 197684 343272 197736
rect 343324 197724 343330 197736
rect 343450 197724 343456 197736
rect 343324 197696 343456 197724
rect 343324 197684 343330 197696
rect 343450 197684 343456 197696
rect 343508 197684 343514 197736
rect 348970 197684 348976 197736
rect 349028 197724 349034 197736
rect 358078 197724 358084 197736
rect 349028 197696 358084 197724
rect 349028 197684 349034 197696
rect 358078 197684 358084 197696
rect 358136 197684 358142 197736
rect 359366 197684 359372 197736
rect 359424 197724 359430 197736
rect 371878 197724 371884 197736
rect 359424 197696 371884 197724
rect 359424 197684 359430 197696
rect 371878 197684 371884 197696
rect 371936 197684 371942 197736
rect 376662 197684 376668 197736
rect 376720 197724 376726 197736
rect 378888 197724 378916 197764
rect 397089 197761 397101 197795
rect 397135 197792 397147 197795
rect 400858 197792 400864 197804
rect 397135 197764 400864 197792
rect 397135 197761 397147 197764
rect 397089 197755 397147 197761
rect 400858 197752 400864 197764
rect 400916 197752 400922 197804
rect 402946 197792 402974 197832
rect 403250 197820 403256 197872
rect 403308 197860 403314 197872
rect 472618 197860 472624 197872
rect 403308 197832 472624 197860
rect 403308 197820 403314 197832
rect 472618 197820 472624 197832
rect 472676 197820 472682 197872
rect 407761 197795 407819 197801
rect 407761 197792 407773 197795
rect 402946 197764 407773 197792
rect 407761 197761 407773 197764
rect 407807 197761 407819 197795
rect 407761 197755 407819 197761
rect 409506 197752 409512 197804
rect 409564 197792 409570 197804
rect 478138 197792 478144 197804
rect 409564 197764 478144 197792
rect 409564 197752 409570 197764
rect 478138 197752 478144 197764
rect 478196 197752 478202 197804
rect 376720 197696 378916 197724
rect 376720 197684 376726 197696
rect 380066 197684 380072 197736
rect 380124 197724 380130 197736
rect 380124 197696 404768 197724
rect 380124 197684 380130 197696
rect 98638 197616 98644 197668
rect 98696 197656 98702 197668
rect 198182 197656 198188 197668
rect 98696 197628 198188 197656
rect 98696 197616 98702 197628
rect 198182 197616 198188 197628
rect 198240 197616 198246 197668
rect 199378 197616 199384 197668
rect 199436 197656 199442 197668
rect 211614 197656 211620 197668
rect 199436 197628 211620 197656
rect 199436 197616 199442 197628
rect 211614 197616 211620 197628
rect 211672 197616 211678 197668
rect 213178 197616 213184 197668
rect 213236 197656 213242 197668
rect 235994 197656 236000 197668
rect 213236 197628 236000 197656
rect 213236 197616 213242 197628
rect 235994 197616 236000 197628
rect 236052 197616 236058 197668
rect 246298 197616 246304 197668
rect 246356 197656 246362 197668
rect 259638 197656 259644 197668
rect 246356 197628 259644 197656
rect 246356 197616 246362 197628
rect 259638 197616 259644 197628
rect 259696 197616 259702 197668
rect 260742 197616 260748 197668
rect 260800 197656 260806 197668
rect 279142 197656 279148 197668
rect 260800 197628 279148 197656
rect 260800 197616 260806 197628
rect 279142 197616 279148 197628
rect 279200 197616 279206 197668
rect 358354 197616 358360 197668
rect 358412 197656 358418 197668
rect 364886 197656 364892 197668
rect 358412 197628 364892 197656
rect 358412 197616 358418 197628
rect 364886 197616 364892 197628
rect 364944 197616 364950 197668
rect 365530 197616 365536 197668
rect 365588 197656 365594 197668
rect 372062 197656 372068 197668
rect 365588 197628 372068 197656
rect 365588 197616 365594 197628
rect 372062 197616 372068 197628
rect 372120 197616 372126 197668
rect 372338 197616 372344 197668
rect 372396 197656 372402 197668
rect 381446 197656 381452 197668
rect 372396 197628 381452 197656
rect 372396 197616 372402 197628
rect 381446 197616 381452 197628
rect 381504 197616 381510 197668
rect 383194 197616 383200 197668
rect 383252 197656 383258 197668
rect 404740 197656 404768 197696
rect 405458 197684 405464 197736
rect 405516 197724 405522 197736
rect 405642 197724 405648 197736
rect 405516 197696 405648 197724
rect 405516 197684 405522 197696
rect 405642 197684 405648 197696
rect 405700 197684 405706 197736
rect 412542 197684 412548 197736
rect 412600 197724 412606 197736
rect 479518 197724 479524 197736
rect 412600 197696 479524 197724
rect 412600 197684 412606 197696
rect 479518 197684 479524 197696
rect 479576 197684 479582 197736
rect 406470 197656 406476 197668
rect 383252 197628 402974 197656
rect 404740 197628 406476 197656
rect 383252 197616 383258 197628
rect 105538 197548 105544 197600
rect 105596 197588 105602 197600
rect 201494 197588 201500 197600
rect 105596 197560 201500 197588
rect 105596 197548 105602 197560
rect 201494 197548 201500 197560
rect 201552 197548 201558 197600
rect 215938 197548 215944 197600
rect 215996 197588 216002 197600
rect 222194 197588 222200 197600
rect 215996 197560 222200 197588
rect 215996 197548 216002 197560
rect 222194 197548 222200 197560
rect 222252 197548 222258 197600
rect 224218 197548 224224 197600
rect 224276 197588 224282 197600
rect 243078 197588 243084 197600
rect 224276 197560 243084 197588
rect 224276 197548 224282 197560
rect 243078 197548 243084 197560
rect 243136 197548 243142 197600
rect 263134 197588 263140 197600
rect 258046 197560 263140 197588
rect 125502 197480 125508 197532
rect 125560 197520 125566 197532
rect 219894 197520 219900 197532
rect 125560 197492 219900 197520
rect 125560 197480 125566 197492
rect 219894 197480 219900 197492
rect 219952 197480 219958 197532
rect 256050 197480 256056 197532
rect 256108 197520 256114 197532
rect 258046 197520 258074 197560
rect 263134 197548 263140 197560
rect 263192 197548 263198 197600
rect 267090 197548 267096 197600
rect 267148 197588 267154 197600
rect 271414 197588 271420 197600
rect 267148 197560 271420 197588
rect 267148 197548 267154 197560
rect 271414 197548 271420 197560
rect 271472 197548 271478 197600
rect 300762 197548 300768 197600
rect 300820 197588 300826 197600
rect 305638 197588 305644 197600
rect 300820 197560 305644 197588
rect 300820 197548 300826 197560
rect 305638 197548 305644 197560
rect 305696 197548 305702 197600
rect 309042 197548 309048 197600
rect 309100 197588 309106 197600
rect 309870 197588 309876 197600
rect 309100 197560 309876 197588
rect 309100 197548 309106 197560
rect 309870 197548 309876 197560
rect 309928 197548 309934 197600
rect 312354 197548 312360 197600
rect 312412 197588 312418 197600
rect 313918 197588 313924 197600
rect 312412 197560 313924 197588
rect 312412 197548 312418 197560
rect 313918 197548 313924 197560
rect 313976 197548 313982 197600
rect 321094 197548 321100 197600
rect 321152 197588 321158 197600
rect 321370 197588 321376 197600
rect 321152 197560 321376 197588
rect 321152 197548 321158 197560
rect 321370 197548 321376 197560
rect 321428 197548 321434 197600
rect 325418 197548 325424 197600
rect 325476 197588 325482 197600
rect 325602 197588 325608 197600
rect 325476 197560 325608 197588
rect 325476 197548 325482 197560
rect 325602 197548 325608 197560
rect 325660 197548 325666 197600
rect 364150 197548 364156 197600
rect 364208 197588 364214 197600
rect 376018 197588 376024 197600
rect 364208 197560 376024 197588
rect 364208 197548 364214 197560
rect 376018 197548 376024 197560
rect 376076 197548 376082 197600
rect 384666 197548 384672 197600
rect 384724 197588 384730 197600
rect 388438 197588 388444 197600
rect 384724 197560 388444 197588
rect 384724 197548 384730 197560
rect 388438 197548 388444 197560
rect 388496 197548 388502 197600
rect 394881 197591 394939 197597
rect 388548 197560 394832 197588
rect 256108 197492 258074 197520
rect 256108 197480 256114 197492
rect 260098 197480 260104 197532
rect 260156 197520 260162 197532
rect 269942 197520 269948 197532
rect 260156 197492 267734 197520
rect 260156 197480 260162 197492
rect 111058 197412 111064 197464
rect 111116 197452 111122 197464
rect 111116 197424 200114 197452
rect 111116 197412 111122 197424
rect 173158 197344 173164 197396
rect 173216 197384 173222 197396
rect 177574 197384 177580 197396
rect 173216 197356 177580 197384
rect 173216 197344 173222 197356
rect 177574 197344 177580 197356
rect 177632 197344 177638 197396
rect 181438 197344 181444 197396
rect 181496 197384 181502 197396
rect 185302 197384 185308 197396
rect 181496 197356 185308 197384
rect 181496 197344 181502 197356
rect 185302 197344 185308 197356
rect 185360 197344 185366 197396
rect 186958 197344 186964 197396
rect 187016 197384 187022 197396
rect 199654 197384 199660 197396
rect 187016 197356 199660 197384
rect 187016 197344 187022 197356
rect 199654 197344 199660 197356
rect 199712 197344 199718 197396
rect 200086 197384 200114 197424
rect 202138 197412 202144 197464
rect 202196 197452 202202 197464
rect 208486 197452 208492 197464
rect 202196 197424 208492 197452
rect 202196 197412 202202 197424
rect 208486 197412 208492 197424
rect 208544 197412 208550 197464
rect 264238 197412 264244 197464
rect 264296 197452 264302 197464
rect 265710 197452 265716 197464
rect 264296 197424 265716 197452
rect 264296 197412 264302 197424
rect 265710 197412 265716 197424
rect 265768 197412 265774 197464
rect 267706 197452 267734 197492
rect 268120 197492 269948 197520
rect 268120 197452 268148 197492
rect 269942 197480 269948 197492
rect 270000 197480 270006 197532
rect 296346 197480 296352 197532
rect 296404 197520 296410 197532
rect 298094 197520 298100 197532
rect 296404 197492 298100 197520
rect 296404 197480 296410 197492
rect 298094 197480 298100 197492
rect 298152 197480 298158 197532
rect 302050 197480 302056 197532
rect 302108 197520 302114 197532
rect 304258 197520 304264 197532
rect 302108 197492 304264 197520
rect 302108 197480 302114 197492
rect 304258 197480 304264 197492
rect 304316 197480 304322 197532
rect 315482 197480 315488 197532
rect 315540 197520 315546 197532
rect 318150 197520 318156 197532
rect 315540 197492 318156 197520
rect 315540 197480 315546 197492
rect 318150 197480 318156 197492
rect 318208 197480 318214 197532
rect 324222 197480 324228 197532
rect 324280 197520 324286 197532
rect 356698 197520 356704 197532
rect 324280 197492 356704 197520
rect 324280 197480 324286 197492
rect 356698 197480 356704 197492
rect 356756 197480 356762 197532
rect 358814 197480 358820 197532
rect 358872 197520 358878 197532
rect 359550 197520 359556 197532
rect 358872 197492 359556 197520
rect 358872 197480 358878 197492
rect 359550 197480 359556 197492
rect 359608 197480 359614 197532
rect 362402 197480 362408 197532
rect 362460 197520 362466 197532
rect 366358 197520 366364 197532
rect 362460 197492 366364 197520
rect 362460 197480 362466 197492
rect 366358 197480 366364 197492
rect 366416 197480 366422 197532
rect 371786 197480 371792 197532
rect 371844 197520 371850 197532
rect 385678 197520 385684 197532
rect 371844 197492 385684 197520
rect 371844 197480 371850 197492
rect 385678 197480 385684 197492
rect 385736 197480 385742 197532
rect 386138 197480 386144 197532
rect 386196 197520 386202 197532
rect 388548 197520 388576 197560
rect 386196 197492 388576 197520
rect 386196 197480 386202 197492
rect 389082 197480 389088 197532
rect 389140 197520 389146 197532
rect 394804 197520 394832 197560
rect 394881 197557 394893 197591
rect 394927 197588 394939 197591
rect 396718 197588 396724 197600
rect 394927 197560 396724 197588
rect 394927 197557 394939 197560
rect 394881 197551 394939 197557
rect 396718 197548 396724 197560
rect 396776 197548 396782 197600
rect 399202 197548 399208 197600
rect 399260 197588 399266 197600
rect 400122 197588 400128 197600
rect 399260 197560 400128 197588
rect 399260 197548 399266 197560
rect 400122 197548 400128 197560
rect 400180 197548 400186 197600
rect 402946 197588 402974 197628
rect 406470 197616 406476 197628
rect 406528 197616 406534 197668
rect 406562 197616 406568 197668
rect 406620 197656 406626 197668
rect 406620 197628 412634 197656
rect 406620 197616 406626 197628
rect 407758 197588 407764 197600
rect 402946 197560 407764 197588
rect 407758 197548 407764 197560
rect 407816 197548 407822 197600
rect 407850 197548 407856 197600
rect 407908 197588 407914 197600
rect 409138 197588 409144 197600
rect 407908 197560 409144 197588
rect 407908 197548 407914 197560
rect 409138 197548 409144 197560
rect 409196 197548 409202 197600
rect 410886 197548 410892 197600
rect 410944 197588 410950 197600
rect 411162 197588 411168 197600
rect 410944 197560 411168 197588
rect 410944 197548 410950 197560
rect 411162 197548 411168 197560
rect 411220 197548 411226 197600
rect 412606 197588 412634 197628
rect 415302 197616 415308 197668
rect 415360 197656 415366 197668
rect 415360 197628 423076 197656
rect 415360 197616 415366 197628
rect 412606 197560 422892 197588
rect 397089 197523 397147 197529
rect 397089 197520 397101 197523
rect 389140 197492 393314 197520
rect 394804 197492 397101 197520
rect 389140 197480 389146 197492
rect 267706 197424 268148 197452
rect 269758 197412 269764 197464
rect 269816 197452 269822 197464
rect 271966 197452 271972 197464
rect 269816 197424 271972 197452
rect 269816 197412 269822 197424
rect 271966 197412 271972 197424
rect 272024 197412 272030 197464
rect 282178 197412 282184 197464
rect 282236 197452 282242 197464
rect 284846 197452 284852 197464
rect 282236 197424 284852 197452
rect 282236 197412 282242 197424
rect 284846 197412 284852 197424
rect 284904 197412 284910 197464
rect 284938 197412 284944 197464
rect 284996 197452 285002 197464
rect 286502 197452 286508 197464
rect 284996 197424 286508 197452
rect 284996 197412 285002 197424
rect 286502 197412 286508 197424
rect 286560 197412 286566 197464
rect 300026 197412 300032 197464
rect 300084 197452 300090 197464
rect 300762 197452 300768 197464
rect 300084 197424 300768 197452
rect 300084 197412 300090 197424
rect 300762 197412 300768 197424
rect 300820 197412 300826 197464
rect 301498 197412 301504 197464
rect 301556 197452 301562 197464
rect 307018 197452 307024 197464
rect 301556 197424 307024 197452
rect 301556 197412 301562 197424
rect 307018 197412 307024 197424
rect 307076 197412 307082 197464
rect 314930 197412 314936 197464
rect 314988 197452 314994 197464
rect 316678 197452 316684 197464
rect 314988 197424 316684 197452
rect 314988 197412 314994 197424
rect 316678 197412 316684 197424
rect 316736 197412 316742 197464
rect 323210 197412 323216 197464
rect 323268 197452 323274 197464
rect 324130 197452 324136 197464
rect 323268 197424 324136 197452
rect 323268 197412 323274 197424
rect 324130 197412 324136 197424
rect 324188 197412 324194 197464
rect 332042 197412 332048 197464
rect 332100 197452 332106 197464
rect 332502 197452 332508 197464
rect 332100 197424 332508 197452
rect 332100 197412 332106 197424
rect 332502 197412 332508 197424
rect 332560 197412 332566 197464
rect 334618 197412 334624 197464
rect 334676 197452 334682 197464
rect 335170 197452 335176 197464
rect 334676 197424 335176 197452
rect 334676 197412 334682 197424
rect 335170 197412 335176 197424
rect 335228 197412 335234 197464
rect 336090 197412 336096 197464
rect 336148 197452 336154 197464
rect 341610 197452 341616 197464
rect 336148 197424 341616 197452
rect 336148 197412 336154 197424
rect 341610 197412 341616 197424
rect 341668 197412 341674 197464
rect 345474 197412 345480 197464
rect 345532 197452 345538 197464
rect 346210 197452 346216 197464
rect 345532 197424 346216 197452
rect 345532 197412 345538 197424
rect 346210 197412 346216 197424
rect 346268 197412 346274 197464
rect 351178 197412 351184 197464
rect 351236 197452 351242 197464
rect 356790 197452 356796 197464
rect 351236 197424 356796 197452
rect 351236 197412 351242 197424
rect 356790 197412 356796 197424
rect 356848 197412 356854 197464
rect 361482 197412 361488 197464
rect 361540 197452 361546 197464
rect 363598 197452 363604 197464
rect 361540 197424 363604 197452
rect 361540 197412 361546 197424
rect 363598 197412 363604 197424
rect 363656 197412 363662 197464
rect 364058 197412 364064 197464
rect 364116 197452 364122 197464
rect 370682 197452 370688 197464
rect 364116 197424 370688 197452
rect 364116 197412 364122 197424
rect 370682 197412 370688 197424
rect 370740 197412 370746 197464
rect 373258 197412 373264 197464
rect 373316 197452 373322 197464
rect 374638 197452 374644 197464
rect 373316 197424 374644 197452
rect 373316 197412 373322 197424
rect 374638 197412 374644 197424
rect 374696 197412 374702 197464
rect 374914 197412 374920 197464
rect 374972 197452 374978 197464
rect 377398 197452 377404 197464
rect 374972 197424 377404 197452
rect 374972 197412 374978 197424
rect 377398 197412 377404 197424
rect 377456 197412 377462 197464
rect 387702 197412 387708 197464
rect 387760 197452 387766 197464
rect 388530 197452 388536 197464
rect 387760 197424 388536 197452
rect 387760 197412 387766 197424
rect 388530 197412 388536 197424
rect 388588 197412 388594 197464
rect 389818 197412 389824 197464
rect 389876 197452 389882 197464
rect 390462 197452 390468 197464
rect 389876 197424 390468 197452
rect 389876 197412 389882 197424
rect 390462 197412 390468 197424
rect 390520 197412 390526 197464
rect 393286 197452 393314 197492
rect 397089 197489 397101 197492
rect 397135 197489 397147 197523
rect 397089 197483 397147 197489
rect 398650 197480 398656 197532
rect 398708 197520 398714 197532
rect 399478 197520 399484 197532
rect 398708 197492 399484 197520
rect 398708 197480 398714 197492
rect 399478 197480 399484 197492
rect 399536 197480 399542 197532
rect 399588 197492 401640 197520
rect 399588 197452 399616 197492
rect 401612 197452 401640 197492
rect 402146 197480 402152 197532
rect 402204 197520 402210 197532
rect 402882 197520 402888 197532
rect 402204 197492 402888 197520
rect 402204 197480 402210 197492
rect 402882 197480 402888 197492
rect 402940 197480 402946 197532
rect 403802 197480 403808 197532
rect 403860 197520 403866 197532
rect 404262 197520 404268 197532
rect 403860 197492 404268 197520
rect 403860 197480 403866 197492
rect 404262 197480 404268 197492
rect 404320 197480 404326 197532
rect 404906 197480 404912 197532
rect 404964 197520 404970 197532
rect 406378 197520 406384 197532
rect 404964 197492 406384 197520
rect 404964 197480 404970 197492
rect 406378 197480 406384 197492
rect 406436 197480 406442 197532
rect 407482 197480 407488 197532
rect 407540 197520 407546 197532
rect 408310 197520 408316 197532
rect 407540 197492 408316 197520
rect 407540 197480 407546 197492
rect 408310 197480 408316 197492
rect 408368 197480 408374 197532
rect 408954 197480 408960 197532
rect 409012 197520 409018 197532
rect 409690 197520 409696 197532
rect 409012 197492 409696 197520
rect 409012 197480 409018 197492
rect 409690 197480 409696 197492
rect 409748 197480 409754 197532
rect 410426 197480 410432 197532
rect 410484 197520 410490 197532
rect 410978 197520 410984 197532
rect 410484 197492 410984 197520
rect 410484 197480 410490 197492
rect 410978 197480 410984 197492
rect 411036 197480 411042 197532
rect 412082 197480 412088 197532
rect 412140 197520 412146 197532
rect 412542 197520 412548 197532
rect 412140 197492 412548 197520
rect 412140 197480 412146 197492
rect 412542 197480 412548 197492
rect 412600 197480 412606 197532
rect 418890 197520 418896 197532
rect 412836 197492 418896 197520
rect 412836 197452 412864 197492
rect 418890 197480 418896 197492
rect 418948 197480 418954 197532
rect 420181 197523 420239 197529
rect 420181 197489 420193 197523
rect 420227 197520 420239 197523
rect 422294 197520 422300 197532
rect 420227 197492 422300 197520
rect 420227 197489 420239 197492
rect 420181 197483 420239 197489
rect 422294 197480 422300 197492
rect 422352 197480 422358 197532
rect 393286 197424 399616 197452
rect 400324 197424 401548 197452
rect 401612 197424 412864 197452
rect 412928 197424 416820 197452
rect 202966 197384 202972 197396
rect 200086 197356 202972 197384
rect 202966 197344 202972 197356
rect 203024 197344 203030 197396
rect 204898 197344 204904 197396
rect 204956 197384 204962 197396
rect 205634 197384 205640 197396
rect 204956 197356 205640 197384
rect 204956 197344 204962 197356
rect 205634 197344 205640 197356
rect 205692 197344 205698 197396
rect 206278 197344 206284 197396
rect 206336 197384 206342 197396
rect 207014 197384 207020 197396
rect 206336 197356 207020 197384
rect 206336 197344 206342 197356
rect 207014 197344 207020 197356
rect 207072 197344 207078 197396
rect 220170 197344 220176 197396
rect 220228 197384 220234 197396
rect 223942 197384 223948 197396
rect 220228 197356 223948 197384
rect 220228 197344 220234 197356
rect 223942 197344 223948 197356
rect 224000 197344 224006 197396
rect 244918 197344 244924 197396
rect 244976 197384 244982 197396
rect 247678 197384 247684 197396
rect 244976 197356 247684 197384
rect 244976 197344 244982 197356
rect 247678 197344 247684 197356
rect 247736 197344 247742 197396
rect 250438 197344 250444 197396
rect 250496 197384 250502 197396
rect 253934 197384 253940 197396
rect 250496 197356 253940 197384
rect 250496 197344 250502 197356
rect 253934 197344 253940 197356
rect 253992 197344 253998 197396
rect 262858 197344 262864 197396
rect 262916 197384 262922 197396
rect 264330 197384 264336 197396
rect 262916 197356 264336 197384
rect 262916 197344 262922 197356
rect 264330 197344 264336 197356
rect 264388 197344 264394 197396
rect 266998 197344 267004 197396
rect 267056 197384 267062 197396
rect 269114 197384 269120 197396
rect 267056 197356 269120 197384
rect 267056 197344 267062 197356
rect 269114 197344 269120 197356
rect 269172 197344 269178 197396
rect 269850 197344 269856 197396
rect 269908 197384 269914 197396
rect 270862 197384 270868 197396
rect 269908 197356 270868 197384
rect 269908 197344 269914 197356
rect 270862 197344 270868 197356
rect 270920 197344 270926 197396
rect 271138 197344 271144 197396
rect 271196 197384 271202 197396
rect 273622 197384 273628 197396
rect 271196 197356 273628 197384
rect 271196 197344 271202 197356
rect 273622 197344 273628 197356
rect 273680 197344 273686 197396
rect 273898 197344 273904 197396
rect 273956 197384 273962 197396
rect 275094 197384 275100 197396
rect 273956 197356 275100 197384
rect 273956 197344 273962 197356
rect 275094 197344 275100 197356
rect 275152 197344 275158 197396
rect 280798 197344 280804 197396
rect 280856 197384 280862 197396
rect 281534 197384 281540 197396
rect 280856 197356 281540 197384
rect 280856 197344 280862 197356
rect 281534 197344 281540 197356
rect 281592 197344 281598 197396
rect 282270 197344 282276 197396
rect 282328 197384 282334 197396
rect 284294 197384 284300 197396
rect 282328 197356 284300 197384
rect 282328 197344 282334 197356
rect 284294 197344 284300 197356
rect 284352 197344 284358 197396
rect 286318 197344 286324 197396
rect 286376 197384 286382 197396
rect 287422 197384 287428 197396
rect 286376 197356 287428 197384
rect 286376 197344 286382 197356
rect 287422 197344 287428 197356
rect 287480 197344 287486 197396
rect 287698 197344 287704 197396
rect 287756 197384 287762 197396
rect 289078 197384 289084 197396
rect 287756 197356 289084 197384
rect 287756 197344 287762 197356
rect 289078 197344 289084 197356
rect 289136 197344 289142 197396
rect 289722 197344 289728 197396
rect 289780 197384 289786 197396
rect 291654 197384 291660 197396
rect 289780 197356 291660 197384
rect 289780 197344 289786 197356
rect 291654 197344 291660 197356
rect 291712 197344 291718 197396
rect 297450 197344 297456 197396
rect 297508 197384 297514 197396
rect 298830 197384 298836 197396
rect 297508 197356 298836 197384
rect 297508 197344 297514 197356
rect 298830 197344 298836 197356
rect 298888 197344 298894 197396
rect 298922 197344 298928 197396
rect 298980 197384 298986 197396
rect 300118 197384 300124 197396
rect 298980 197356 300124 197384
rect 298980 197344 298986 197356
rect 300118 197344 300124 197356
rect 300176 197344 300182 197396
rect 305730 197344 305736 197396
rect 305788 197384 305794 197396
rect 306190 197384 306196 197396
rect 305788 197356 306196 197384
rect 305788 197344 305794 197356
rect 306190 197344 306196 197356
rect 306248 197344 306254 197396
rect 308306 197344 308312 197396
rect 308364 197384 308370 197396
rect 309778 197384 309784 197396
rect 308364 197356 309784 197384
rect 308364 197344 308370 197356
rect 309778 197344 309784 197356
rect 309836 197344 309842 197396
rect 316586 197344 316592 197396
rect 316644 197384 316650 197396
rect 317322 197384 317328 197396
rect 316644 197356 317328 197384
rect 316644 197344 316650 197356
rect 317322 197344 317328 197356
rect 317380 197344 317386 197396
rect 317966 197344 317972 197396
rect 318024 197384 318030 197396
rect 318702 197384 318708 197396
rect 318024 197356 318708 197384
rect 318024 197344 318030 197356
rect 318702 197344 318708 197356
rect 318760 197344 318766 197396
rect 319530 197344 319536 197396
rect 319588 197384 319594 197396
rect 322198 197384 322204 197396
rect 319588 197356 322204 197384
rect 319588 197344 319594 197356
rect 322198 197344 322204 197356
rect 322256 197344 322262 197396
rect 323762 197344 323768 197396
rect 323820 197384 323826 197396
rect 324222 197384 324228 197396
rect 323820 197356 324228 197384
rect 323820 197344 323826 197356
rect 324222 197344 324228 197356
rect 324280 197344 324286 197396
rect 324866 197344 324872 197396
rect 324924 197384 324930 197396
rect 325418 197384 325424 197396
rect 324924 197356 325424 197384
rect 324924 197344 324930 197356
rect 325418 197344 325424 197356
rect 325476 197344 325482 197396
rect 327810 197344 327816 197396
rect 327868 197384 327874 197396
rect 328362 197384 328368 197396
rect 327868 197356 328368 197384
rect 327868 197344 327874 197356
rect 328362 197344 328368 197356
rect 328420 197344 328426 197396
rect 330386 197344 330392 197396
rect 330444 197384 330450 197396
rect 331122 197384 331128 197396
rect 330444 197356 331128 197384
rect 330444 197344 330450 197356
rect 331122 197344 331128 197356
rect 331180 197344 331186 197396
rect 331490 197344 331496 197396
rect 331548 197384 331554 197396
rect 332318 197384 332324 197396
rect 331548 197356 332324 197384
rect 331548 197344 331554 197356
rect 332318 197344 332324 197356
rect 332376 197344 332382 197396
rect 334986 197344 334992 197396
rect 335044 197384 335050 197396
rect 335262 197384 335268 197396
rect 335044 197356 335268 197384
rect 335044 197344 335050 197356
rect 335262 197344 335268 197356
rect 335320 197344 335326 197396
rect 337194 197344 337200 197396
rect 337252 197384 337258 197396
rect 338022 197384 338028 197396
rect 337252 197356 338028 197384
rect 337252 197344 337258 197356
rect 338022 197344 338028 197356
rect 338080 197344 338086 197396
rect 338666 197344 338672 197396
rect 338724 197384 338730 197396
rect 339310 197384 339316 197396
rect 338724 197356 339316 197384
rect 338724 197344 338730 197356
rect 339310 197344 339316 197356
rect 339368 197344 339374 197396
rect 341242 197344 341248 197396
rect 341300 197384 341306 197396
rect 342162 197384 342168 197396
rect 341300 197356 342168 197384
rect 341300 197344 341306 197356
rect 342162 197344 342168 197356
rect 342220 197344 342226 197396
rect 342898 197344 342904 197396
rect 342956 197384 342962 197396
rect 343542 197384 343548 197396
rect 342956 197356 343548 197384
rect 342956 197344 342962 197356
rect 343542 197344 343548 197356
rect 343600 197344 343606 197396
rect 346026 197344 346032 197396
rect 346084 197384 346090 197396
rect 346302 197384 346308 197396
rect 346084 197356 346308 197384
rect 346084 197344 346090 197356
rect 346302 197344 346308 197356
rect 346360 197344 346366 197396
rect 346946 197344 346952 197396
rect 347004 197384 347010 197396
rect 347590 197384 347596 197396
rect 347004 197356 347596 197384
rect 347004 197344 347010 197356
rect 347590 197344 347596 197356
rect 347648 197344 347654 197396
rect 348602 197344 348608 197396
rect 348660 197384 348666 197396
rect 349062 197384 349068 197396
rect 348660 197356 349068 197384
rect 348660 197344 348666 197356
rect 349062 197344 349068 197356
rect 349120 197344 349126 197396
rect 349522 197344 349528 197396
rect 349580 197384 349586 197396
rect 350350 197384 350356 197396
rect 349580 197356 350356 197384
rect 349580 197344 349586 197356
rect 350350 197344 350356 197356
rect 350408 197344 350414 197396
rect 352650 197344 352656 197396
rect 352708 197384 352714 197396
rect 353110 197384 353116 197396
rect 352708 197356 353116 197384
rect 352708 197344 352714 197356
rect 353110 197344 353116 197356
rect 353168 197344 353174 197396
rect 355226 197344 355232 197396
rect 355284 197384 355290 197396
rect 360838 197384 360844 197396
rect 355284 197356 360844 197384
rect 355284 197344 355290 197356
rect 360838 197344 360844 197356
rect 360896 197344 360902 197396
rect 362034 197344 362040 197396
rect 362092 197384 362098 197396
rect 362862 197384 362868 197396
rect 362092 197356 362868 197384
rect 362092 197344 362098 197356
rect 362862 197344 362868 197356
rect 362920 197344 362926 197396
rect 363506 197344 363512 197396
rect 363564 197384 363570 197396
rect 364242 197384 364248 197396
rect 363564 197356 364248 197384
rect 363564 197344 363570 197356
rect 364242 197344 364248 197356
rect 364300 197344 364306 197396
rect 364978 197344 364984 197396
rect 365036 197384 365042 197396
rect 365622 197384 365628 197396
rect 365036 197356 365628 197384
rect 365036 197344 365042 197356
rect 365622 197344 365628 197356
rect 365680 197344 365686 197396
rect 368382 197344 368388 197396
rect 368440 197384 368446 197396
rect 370498 197384 370504 197396
rect 368440 197356 370504 197384
rect 368440 197344 368446 197356
rect 370498 197344 370504 197356
rect 370556 197344 370562 197396
rect 374362 197344 374368 197396
rect 374420 197384 374426 197396
rect 375190 197384 375196 197396
rect 374420 197356 375196 197384
rect 374420 197344 374426 197356
rect 375190 197344 375196 197356
rect 375248 197344 375254 197396
rect 375834 197344 375840 197396
rect 375892 197384 375898 197396
rect 376386 197384 376392 197396
rect 375892 197356 376392 197384
rect 375892 197344 375898 197356
rect 376386 197344 376392 197356
rect 376444 197344 376450 197396
rect 377490 197344 377496 197396
rect 377548 197384 377554 197396
rect 377950 197384 377956 197396
rect 377548 197356 377956 197384
rect 377548 197344 377554 197356
rect 377950 197344 377956 197356
rect 378008 197344 378014 197396
rect 378410 197344 378416 197396
rect 378468 197384 378474 197396
rect 379238 197384 379244 197396
rect 378468 197356 379244 197384
rect 378468 197344 378474 197356
rect 379238 197344 379244 197356
rect 379296 197344 379302 197396
rect 381538 197344 381544 197396
rect 381596 197384 381602 197396
rect 382090 197384 382096 197396
rect 381596 197356 382096 197384
rect 381596 197344 381602 197356
rect 382090 197344 382096 197356
rect 382148 197344 382154 197396
rect 382642 197344 382648 197396
rect 382700 197384 382706 197396
rect 383562 197384 383568 197396
rect 382700 197356 383568 197384
rect 382700 197344 382706 197356
rect 383562 197344 383568 197356
rect 383620 197344 383626 197396
rect 384114 197344 384120 197396
rect 384172 197384 384178 197396
rect 384942 197384 384948 197396
rect 384172 197356 384948 197384
rect 384172 197344 384178 197356
rect 384942 197344 384948 197356
rect 385000 197344 385006 197396
rect 385770 197344 385776 197396
rect 385828 197384 385834 197396
rect 386322 197384 386328 197396
rect 385828 197356 386328 197384
rect 385828 197344 385834 197356
rect 386322 197344 386328 197356
rect 386380 197344 386386 197396
rect 388346 197344 388352 197396
rect 388404 197384 388410 197396
rect 388806 197384 388812 197396
rect 388404 197356 388812 197384
rect 388404 197344 388410 197356
rect 388806 197344 388812 197356
rect 388864 197344 388870 197396
rect 390922 197344 390928 197396
rect 390980 197384 390986 197396
rect 392578 197384 392584 197396
rect 390980 197356 392584 197384
rect 390980 197344 390986 197356
rect 392578 197344 392584 197356
rect 392636 197344 392642 197396
rect 393038 197344 393044 197396
rect 393096 197384 393102 197396
rect 393222 197384 393228 197396
rect 393096 197356 393228 197384
rect 393096 197344 393102 197356
rect 393222 197344 393228 197356
rect 393280 197344 393286 197396
rect 394050 197344 394056 197396
rect 394108 197384 394114 197396
rect 395338 197384 395344 197396
rect 394108 197356 395344 197384
rect 394108 197344 394114 197356
rect 395338 197344 395344 197356
rect 395396 197344 395402 197396
rect 396626 197344 396632 197396
rect 396684 197384 396690 197396
rect 397270 197384 397276 197396
rect 396684 197356 397276 197384
rect 396684 197344 396690 197356
rect 397270 197344 397276 197356
rect 397328 197344 397334 197396
rect 398098 197344 398104 197396
rect 398156 197384 398162 197396
rect 398742 197384 398748 197396
rect 398156 197356 398748 197384
rect 398156 197344 398162 197356
rect 398742 197344 398748 197356
rect 398800 197344 398806 197396
rect 399570 197344 399576 197396
rect 399628 197384 399634 197396
rect 400030 197384 400036 197396
rect 399628 197356 400036 197384
rect 399628 197344 399634 197356
rect 400030 197344 400036 197356
rect 400088 197344 400094 197396
rect 400125 197387 400183 197393
rect 400125 197353 400137 197387
rect 400171 197384 400183 197387
rect 400324 197384 400352 197424
rect 400171 197356 400352 197384
rect 400171 197353 400183 197356
rect 400125 197347 400183 197353
rect 400674 197344 400680 197396
rect 400732 197384 400738 197396
rect 401410 197384 401416 197396
rect 400732 197356 401416 197384
rect 400732 197344 400738 197356
rect 401410 197344 401416 197356
rect 401468 197344 401474 197396
rect 401520 197384 401548 197424
rect 412928 197384 412956 197424
rect 401520 197356 412956 197384
rect 413002 197344 413008 197396
rect 413060 197384 413066 197396
rect 413830 197384 413836 197396
rect 413060 197356 413836 197384
rect 413060 197344 413066 197356
rect 413830 197344 413836 197356
rect 413888 197344 413894 197396
rect 414658 197344 414664 197396
rect 414716 197384 414722 197396
rect 415302 197384 415308 197396
rect 414716 197356 415308 197384
rect 414716 197344 414722 197356
rect 415302 197344 415308 197356
rect 415360 197344 415366 197396
rect 416130 197344 416136 197396
rect 416188 197384 416194 197396
rect 416682 197384 416688 197396
rect 416188 197356 416688 197384
rect 416188 197344 416194 197356
rect 416682 197344 416688 197356
rect 416740 197344 416746 197396
rect 416792 197384 416820 197424
rect 417234 197412 417240 197464
rect 417292 197452 417298 197464
rect 418798 197452 418804 197464
rect 417292 197424 418804 197452
rect 417292 197412 417298 197424
rect 418798 197412 418804 197424
rect 418856 197412 418862 197464
rect 422864 197452 422892 197560
rect 423048 197520 423076 197628
rect 428645 197591 428703 197597
rect 428645 197557 428657 197591
rect 428691 197588 428703 197591
rect 473998 197588 474004 197600
rect 428691 197560 474004 197588
rect 428691 197557 428703 197560
rect 428645 197551 428703 197557
rect 473998 197548 474004 197560
rect 474056 197548 474062 197600
rect 482278 197520 482284 197532
rect 423048 197492 429884 197520
rect 428645 197455 428703 197461
rect 428645 197452 428657 197455
rect 422864 197424 428657 197452
rect 428645 197421 428657 197424
rect 428691 197421 428703 197455
rect 429856 197452 429884 197492
rect 434686 197492 482284 197520
rect 434686 197452 434714 197492
rect 482278 197480 482284 197492
rect 482336 197480 482342 197532
rect 429856 197424 434714 197452
rect 428645 197415 428703 197421
rect 417418 197384 417424 197396
rect 416792 197356 417424 197384
rect 417418 197344 417424 197356
rect 417476 197344 417482 197396
rect 417786 197344 417792 197396
rect 417844 197384 417850 197396
rect 418062 197384 418068 197396
rect 417844 197356 418068 197384
rect 417844 197344 417850 197356
rect 418062 197344 418068 197356
rect 418120 197344 418126 197396
rect 418706 197344 418712 197396
rect 418764 197384 418770 197396
rect 486418 197384 486424 197396
rect 418764 197356 486424 197384
rect 418764 197344 418770 197356
rect 486418 197344 486424 197356
rect 486476 197344 486482 197396
rect 200758 196868 200764 196920
rect 200816 196908 200822 196920
rect 242986 196908 242992 196920
rect 200816 196880 242992 196908
rect 200816 196868 200822 196880
rect 242986 196868 242992 196880
rect 243044 196868 243050 196920
rect 169570 196800 169576 196852
rect 169628 196840 169634 196852
rect 238938 196840 238944 196852
rect 169628 196812 238944 196840
rect 169628 196800 169634 196812
rect 238938 196800 238944 196812
rect 238996 196800 239002 196852
rect 88242 196732 88248 196784
rect 88300 196772 88306 196784
rect 203886 196772 203892 196784
rect 88300 196744 203892 196772
rect 88300 196732 88306 196744
rect 203886 196732 203892 196744
rect 203944 196732 203950 196784
rect 380618 196732 380624 196784
rect 380676 196772 380682 196784
rect 489914 196772 489920 196784
rect 380676 196744 489920 196772
rect 380676 196732 380682 196744
rect 489914 196732 489920 196744
rect 489972 196732 489978 196784
rect 39298 196664 39304 196716
rect 39356 196704 39362 196716
rect 182174 196704 182180 196716
rect 39356 196676 182180 196704
rect 39356 196664 39362 196676
rect 182174 196664 182180 196676
rect 182232 196664 182238 196716
rect 188338 196664 188344 196716
rect 188396 196704 188402 196716
rect 247126 196704 247132 196716
rect 188396 196676 247132 196704
rect 188396 196664 188402 196676
rect 247126 196664 247132 196676
rect 247184 196664 247190 196716
rect 386690 196664 386696 196716
rect 386748 196704 386754 196716
rect 505094 196704 505100 196716
rect 386748 196676 505100 196704
rect 386748 196664 386754 196676
rect 505094 196664 505100 196676
rect 505152 196664 505158 196716
rect 14550 196596 14556 196648
rect 14608 196636 14614 196648
rect 171318 196636 171324 196648
rect 14608 196608 171324 196636
rect 14608 196596 14614 196608
rect 171318 196596 171324 196608
rect 171376 196596 171382 196648
rect 180058 196596 180064 196648
rect 180116 196636 180122 196648
rect 243630 196636 243636 196648
rect 180116 196608 243636 196636
rect 180116 196596 180122 196608
rect 243630 196596 243636 196608
rect 243688 196596 243694 196648
rect 391842 196596 391848 196648
rect 391900 196636 391906 196648
rect 516134 196636 516140 196648
rect 391900 196608 516140 196636
rect 391900 196596 391906 196608
rect 516134 196596 516140 196608
rect 516192 196596 516198 196648
rect 165614 195236 165620 195288
rect 165672 195276 165678 195288
rect 166166 195276 166172 195288
rect 165672 195248 166172 195276
rect 165672 195236 165678 195248
rect 166166 195236 166172 195248
rect 166224 195236 166230 195288
rect 172698 195236 172704 195288
rect 172756 195276 172762 195288
rect 173342 195276 173348 195288
rect 172756 195248 173348 195276
rect 172756 195236 172762 195248
rect 173342 195236 173348 195248
rect 173400 195236 173406 195288
rect 178126 195236 178132 195288
rect 178184 195276 178190 195288
rect 179046 195276 179052 195288
rect 178184 195248 179052 195276
rect 178184 195236 178190 195248
rect 179046 195236 179052 195248
rect 179104 195236 179110 195288
rect 182266 195236 182272 195288
rect 182324 195276 182330 195288
rect 183094 195276 183100 195288
rect 182324 195248 183100 195276
rect 182324 195236 182330 195248
rect 183094 195236 183100 195248
rect 183152 195236 183158 195288
rect 186406 195236 186412 195288
rect 186464 195276 186470 195288
rect 186774 195276 186780 195288
rect 186464 195248 186780 195276
rect 186464 195236 186470 195248
rect 186774 195236 186780 195248
rect 186832 195236 186838 195288
rect 237374 195236 237380 195288
rect 237432 195276 237438 195288
rect 237926 195276 237932 195288
rect 237432 195248 237932 195276
rect 237432 195236 237438 195248
rect 237926 195236 237932 195248
rect 237984 195236 237990 195288
rect 251266 195236 251272 195288
rect 251324 195276 251330 195288
rect 251910 195276 251916 195288
rect 251324 195248 251916 195276
rect 251324 195236 251330 195248
rect 251910 195236 251916 195248
rect 251968 195236 251974 195288
rect 254026 195236 254032 195288
rect 254084 195276 254090 195288
rect 254854 195276 254860 195288
rect 254084 195248 254860 195276
rect 254084 195236 254090 195248
rect 254854 195236 254860 195248
rect 254912 195236 254918 195288
rect 190546 195032 190552 195084
rect 190604 195072 190610 195084
rect 191374 195072 191380 195084
rect 190604 195044 191380 195072
rect 190604 195032 190610 195044
rect 191374 195032 191380 195044
rect 191432 195032 191438 195084
rect 245746 194488 245752 194540
rect 245804 194528 245810 194540
rect 246206 194528 246212 194540
rect 245804 194500 246212 194528
rect 245804 194488 245810 194500
rect 246206 194488 246212 194500
rect 246264 194488 246270 194540
rect 244274 193264 244280 193316
rect 244332 193304 244338 193316
rect 244642 193304 244648 193316
rect 244332 193276 244648 193304
rect 244332 193264 244338 193276
rect 244642 193264 244648 193276
rect 244700 193264 244706 193316
rect 428642 193128 428648 193180
rect 428700 193168 428706 193180
rect 580166 193168 580172 193180
rect 428700 193140 580172 193168
rect 428700 193128 428706 193140
rect 580166 193128 580172 193140
rect 580224 193128 580230 193180
rect 168374 191972 168380 192024
rect 168432 192012 168438 192024
rect 169294 192012 169300 192024
rect 168432 191984 169300 192012
rect 168432 191972 168438 191984
rect 169294 191972 169300 191984
rect 169352 191972 169358 192024
rect 198918 191224 198924 191276
rect 198976 191224 198982 191276
rect 198936 191072 198964 191224
rect 231854 191088 231860 191140
rect 231912 191128 231918 191140
rect 232774 191128 232780 191140
rect 231912 191100 232780 191128
rect 231912 191088 231918 191100
rect 232774 191088 232780 191100
rect 232832 191088 232838 191140
rect 198918 191020 198924 191072
rect 198976 191020 198982 191072
rect 244366 190884 244372 190936
rect 244424 190924 244430 190936
rect 245102 190924 245108 190936
rect 244424 190896 245108 190924
rect 244424 190884 244430 190896
rect 245102 190884 245108 190896
rect 245160 190884 245166 190936
rect 2774 188844 2780 188896
rect 2832 188884 2838 188896
rect 4798 188884 4804 188896
rect 2832 188856 4804 188884
rect 2832 188844 2838 188856
rect 4798 188844 4804 188856
rect 4856 188844 4862 188896
rect 198826 188368 198832 188420
rect 198884 188408 198890 188420
rect 199010 188408 199016 188420
rect 198884 188380 199016 188408
rect 198884 188368 198890 188380
rect 199010 188368 199016 188380
rect 199068 188368 199074 188420
rect 209682 177284 209688 177336
rect 209740 177324 209746 177336
rect 256786 177324 256792 177336
rect 209740 177296 256792 177324
rect 209740 177284 209746 177296
rect 256786 177284 256792 177296
rect 256844 177284 256850 177336
rect 258718 176672 258724 176724
rect 258776 176712 258782 176724
rect 266538 176712 266544 176724
rect 258776 176684 266544 176712
rect 258776 176672 258782 176684
rect 266538 176672 266544 176684
rect 266596 176672 266602 176724
rect 220078 171776 220084 171828
rect 220136 171816 220142 171828
rect 258166 171816 258172 171828
rect 220136 171788 258172 171816
rect 220136 171776 220142 171788
rect 258166 171776 258172 171788
rect 258224 171776 258230 171828
rect 424410 166948 424416 167000
rect 424468 166988 424474 167000
rect 580166 166988 580172 167000
rect 424468 166960 580172 166988
rect 424468 166948 424474 166960
rect 580166 166948 580172 166960
rect 580224 166948 580230 167000
rect 3326 164160 3332 164212
rect 3384 164200 3390 164212
rect 10410 164200 10416 164212
rect 3384 164172 10416 164200
rect 3384 164160 3390 164172
rect 10410 164160 10416 164172
rect 10468 164160 10474 164212
rect 204990 155184 204996 155236
rect 205048 155224 205054 155236
rect 244458 155224 244464 155236
rect 205048 155196 244464 155224
rect 205048 155184 205054 155196
rect 244458 155184 244464 155196
rect 244516 155184 244522 155236
rect 428550 153144 428556 153196
rect 428608 153184 428614 153196
rect 580166 153184 580172 153196
rect 428608 153156 580172 153184
rect 428608 153144 428614 153156
rect 580166 153144 580172 153156
rect 580224 153144 580230 153196
rect 3602 150356 3608 150408
rect 3660 150396 3666 150408
rect 100110 150396 100116 150408
rect 3660 150368 100116 150396
rect 3660 150356 3666 150368
rect 100110 150356 100116 150368
rect 100168 150356 100174 150408
rect 429838 139340 429844 139392
rect 429896 139380 429902 139392
rect 580166 139380 580172 139392
rect 429896 139352 580172 139380
rect 429896 139340 429902 139352
rect 580166 139340 580172 139352
rect 580224 139340 580230 139392
rect 421834 126896 421840 126948
rect 421892 126936 421898 126948
rect 580166 126936 580172 126948
rect 421892 126908 580172 126936
rect 421892 126896 421898 126908
rect 580166 126896 580172 126908
rect 580224 126896 580230 126948
rect 425790 113092 425796 113144
rect 425848 113132 425854 113144
rect 579798 113132 579804 113144
rect 425848 113104 579804 113132
rect 425848 113092 425854 113104
rect 579798 113092 579804 113104
rect 579856 113092 579862 113144
rect 3510 110712 3516 110764
rect 3568 110752 3574 110764
rect 7650 110752 7656 110764
rect 3568 110724 7656 110752
rect 3568 110712 3574 110724
rect 7650 110712 7656 110724
rect 7708 110712 7714 110764
rect 428458 100648 428464 100700
rect 428516 100688 428522 100700
rect 580166 100688 580172 100700
rect 428516 100660 580172 100688
rect 428516 100648 428522 100660
rect 580166 100648 580172 100660
rect 580224 100648 580230 100700
rect 3510 97928 3516 97980
rect 3568 97968 3574 97980
rect 101490 97968 101496 97980
rect 3568 97940 101496 97968
rect 3568 97928 3574 97940
rect 101490 97928 101496 97940
rect 101548 97928 101554 97980
rect 103422 89156 103428 89208
rect 103480 89196 103486 89208
rect 210050 89196 210056 89208
rect 103480 89168 210056 89196
rect 103480 89156 103486 89168
rect 210050 89156 210056 89168
rect 210108 89156 210114 89208
rect 81342 89088 81348 89140
rect 81400 89128 81406 89140
rect 200206 89128 200212 89140
rect 81400 89100 200212 89128
rect 81400 89088 81406 89100
rect 200206 89088 200212 89100
rect 200264 89088 200270 89140
rect 35802 89020 35808 89072
rect 35860 89060 35866 89072
rect 170398 89060 170404 89072
rect 35860 89032 170404 89060
rect 35860 89020 35866 89032
rect 170398 89020 170404 89032
rect 170456 89020 170462 89072
rect 23382 88952 23388 89004
rect 23440 88992 23446 89004
rect 175458 88992 175464 89004
rect 23440 88964 175464 88992
rect 23440 88952 23446 88964
rect 175458 88952 175464 88964
rect 175516 88952 175522 89004
rect 384850 88952 384856 89004
rect 384908 88992 384914 89004
rect 500954 88992 500960 89004
rect 384908 88964 500960 88992
rect 384908 88952 384914 88964
rect 500954 88952 500960 88964
rect 501012 88952 501018 89004
rect 135162 87728 135168 87780
rect 135220 87768 135226 87780
rect 220170 87768 220176 87780
rect 135220 87740 220176 87768
rect 135220 87728 135226 87740
rect 220170 87728 220176 87740
rect 220228 87728 220234 87780
rect 43438 87660 43444 87712
rect 43496 87700 43502 87712
rect 183646 87700 183652 87712
rect 43496 87672 183652 87700
rect 43496 87660 43502 87672
rect 183646 87660 183652 87672
rect 183704 87660 183710 87712
rect 28902 87592 28908 87644
rect 28960 87632 28966 87644
rect 173158 87632 173164 87644
rect 28960 87604 173164 87632
rect 28960 87592 28966 87604
rect 173158 87592 173164 87604
rect 173216 87592 173222 87644
rect 242158 87592 242164 87644
rect 242216 87632 242222 87644
rect 265158 87632 265164 87644
rect 242216 87604 265164 87632
rect 242216 87592 242222 87604
rect 265158 87592 265164 87604
rect 265216 87592 265222 87644
rect 372062 87592 372068 87644
rect 372120 87632 372126 87644
rect 456886 87632 456892 87644
rect 372120 87604 456892 87632
rect 372120 87592 372126 87604
rect 456886 87592 456892 87604
rect 456944 87592 456950 87644
rect 421742 86912 421748 86964
rect 421800 86952 421806 86964
rect 580166 86952 580172 86964
rect 421800 86924 580172 86952
rect 421800 86912 421806 86924
rect 580166 86912 580172 86924
rect 580224 86912 580230 86964
rect 341610 86504 341616 86556
rect 341668 86544 341674 86556
rect 389174 86544 389180 86556
rect 341668 86516 389180 86544
rect 341668 86504 341674 86516
rect 389174 86504 389180 86516
rect 389232 86504 389238 86556
rect 366358 86436 366364 86488
rect 366416 86476 366422 86488
rect 448514 86476 448520 86488
rect 366416 86448 448520 86476
rect 366416 86436 366422 86448
rect 448514 86436 448520 86448
rect 448572 86436 448578 86488
rect 362862 86368 362868 86420
rect 362920 86408 362926 86420
rect 448606 86408 448612 86420
rect 362920 86380 448612 86408
rect 362920 86368 362926 86380
rect 448606 86368 448612 86380
rect 448664 86368 448670 86420
rect 379238 86300 379244 86352
rect 379296 86340 379302 86352
rect 485774 86340 485780 86352
rect 379296 86312 485780 86340
rect 379296 86300 379302 86312
rect 485774 86300 485780 86312
rect 485832 86300 485838 86352
rect 106182 86232 106188 86284
rect 106240 86272 106246 86284
rect 199378 86272 199384 86284
rect 106240 86244 199384 86272
rect 106240 86232 106246 86244
rect 199378 86232 199384 86244
rect 199436 86232 199442 86284
rect 206370 86232 206376 86284
rect 206428 86272 206434 86284
rect 252738 86272 252744 86284
rect 206428 86244 252744 86272
rect 206428 86232 206434 86244
rect 252738 86232 252744 86244
rect 252796 86232 252802 86284
rect 340230 86232 340236 86284
rect 340288 86272 340294 86284
rect 382366 86272 382372 86284
rect 340288 86244 382372 86272
rect 340288 86232 340294 86244
rect 382366 86232 382372 86244
rect 382424 86232 382430 86284
rect 388530 86232 388536 86284
rect 388588 86272 388594 86284
rect 506474 86272 506480 86284
rect 388588 86244 506480 86272
rect 388588 86232 388594 86244
rect 506474 86232 506480 86244
rect 506532 86232 506538 86284
rect 3510 85484 3516 85536
rect 3568 85524 3574 85536
rect 64138 85524 64144 85536
rect 3568 85496 64144 85524
rect 3568 85484 3574 85496
rect 64138 85484 64144 85496
rect 64196 85484 64202 85536
rect 162762 85076 162768 85128
rect 162820 85116 162826 85128
rect 216030 85116 216036 85128
rect 162820 85088 216036 85116
rect 162820 85076 162826 85088
rect 216030 85076 216036 85088
rect 216088 85076 216094 85128
rect 143442 85008 143448 85060
rect 143500 85048 143506 85060
rect 217318 85048 217324 85060
rect 143500 85020 217324 85048
rect 143500 85008 143506 85020
rect 217318 85008 217324 85020
rect 217376 85008 217382 85060
rect 113082 84940 113088 84992
rect 113140 84980 113146 84992
rect 197998 84980 198004 84992
rect 113140 84952 198004 84980
rect 113140 84940 113146 84952
rect 197998 84940 198004 84952
rect 198056 84940 198062 84992
rect 198090 84940 198096 84992
rect 198148 84980 198154 84992
rect 251358 84980 251364 84992
rect 198148 84952 251364 84980
rect 198148 84940 198154 84952
rect 251358 84940 251364 84952
rect 251416 84940 251422 84992
rect 137922 84872 137928 84924
rect 137980 84912 137986 84924
rect 225046 84912 225052 84924
rect 137980 84884 225052 84912
rect 137980 84872 137986 84884
rect 225046 84872 225052 84884
rect 225104 84872 225110 84924
rect 370682 84872 370688 84924
rect 370740 84912 370746 84924
rect 452654 84912 452660 84924
rect 370740 84884 452660 84912
rect 370740 84872 370746 84884
rect 452654 84872 452660 84884
rect 452712 84872 452718 84924
rect 95142 84804 95148 84856
rect 95200 84844 95206 84856
rect 206278 84844 206284 84856
rect 95200 84816 206284 84844
rect 95200 84804 95206 84816
rect 206278 84804 206284 84816
rect 206336 84804 206342 84856
rect 400858 84804 400864 84856
rect 400916 84844 400922 84856
rect 503714 84844 503720 84856
rect 400916 84816 503720 84844
rect 400916 84804 400922 84816
rect 503714 84804 503720 84816
rect 503772 84804 503778 84856
rect 147582 80656 147588 80708
rect 147640 80696 147646 80708
rect 213270 80696 213276 80708
rect 147640 80668 213276 80696
rect 147640 80656 147646 80668
rect 213270 80656 213276 80668
rect 213328 80656 213334 80708
rect 424318 73108 424324 73160
rect 424376 73148 424382 73160
rect 580166 73148 580172 73160
rect 424376 73120 580172 73148
rect 424376 73108 424382 73120
rect 580166 73108 580172 73120
rect 580224 73108 580230 73160
rect 3510 71612 3516 71664
rect 3568 71652 3574 71664
rect 7558 71652 7564 71664
rect 3568 71624 7564 71652
rect 3568 71612 3574 71624
rect 7558 71612 7564 71624
rect 7616 71612 7622 71664
rect 425698 60664 425704 60716
rect 425756 60704 425762 60716
rect 580166 60704 580172 60716
rect 425756 60676 580172 60704
rect 425756 60664 425762 60676
rect 580166 60664 580172 60676
rect 580224 60664 580230 60716
rect 3050 59304 3056 59356
rect 3108 59344 3114 59356
rect 100018 59344 100024 59356
rect 3108 59316 100024 59344
rect 3108 59304 3114 59316
rect 100018 59304 100024 59316
rect 100076 59304 100082 59356
rect 421650 46860 421656 46912
rect 421708 46900 421714 46912
rect 580166 46900 580172 46912
rect 421708 46872 580172 46900
rect 421708 46860 421714 46872
rect 580166 46860 580172 46872
rect 580224 46860 580230 46912
rect 3510 45500 3516 45552
rect 3568 45540 3574 45552
rect 82078 45540 82084 45552
rect 3568 45512 82084 45540
rect 3568 45500 3574 45512
rect 82078 45500 82084 45512
rect 82136 45500 82142 45552
rect 99282 44820 99288 44872
rect 99340 44860 99346 44872
rect 202138 44860 202144 44872
rect 99340 44832 202144 44860
rect 99340 44820 99346 44832
rect 202138 44820 202144 44832
rect 202196 44820 202202 44872
rect 385770 44820 385776 44872
rect 385828 44860 385834 44872
rect 470594 44860 470600 44872
rect 385828 44832 470600 44860
rect 385828 44820 385834 44832
rect 470594 44820 470600 44832
rect 470652 44820 470658 44872
rect 370590 35164 370596 35216
rect 370648 35204 370654 35216
rect 438854 35204 438860 35216
rect 370648 35176 438860 35204
rect 370648 35164 370654 35176
rect 438854 35164 438860 35176
rect 438912 35164 438918 35216
rect 2866 33056 2872 33108
rect 2924 33096 2930 33108
rect 10318 33096 10324 33108
rect 2924 33068 10324 33096
rect 2924 33056 2930 33068
rect 10318 33056 10324 33068
rect 10376 33056 10382 33108
rect 508498 33056 508504 33108
rect 508556 33096 508562 33108
rect 580166 33096 580172 33108
rect 508556 33068 580172 33096
rect 508556 33056 508562 33068
rect 580166 33056 580172 33068
rect 580224 33056 580230 33108
rect 388438 26868 388444 26920
rect 388496 26908 388502 26920
rect 499574 26908 499580 26920
rect 388496 26880 499580 26908
rect 388496 26868 388502 26880
rect 499574 26868 499580 26880
rect 499632 26868 499638 26920
rect 370498 25508 370504 25560
rect 370556 25548 370562 25560
rect 463694 25548 463700 25560
rect 370556 25520 463700 25548
rect 370556 25508 370562 25520
rect 463694 25508 463700 25520
rect 463752 25508 463758 25560
rect 392578 24080 392584 24132
rect 392636 24120 392642 24132
rect 514754 24120 514760 24132
rect 392636 24092 514760 24120
rect 392636 24080 392642 24092
rect 514754 24080 514760 24092
rect 514812 24080 514818 24132
rect 245010 22856 245016 22908
rect 245068 22896 245074 22908
rect 267826 22896 267832 22908
rect 245068 22868 267832 22896
rect 245068 22856 245074 22868
rect 267826 22856 267832 22868
rect 267884 22856 267890 22908
rect 216582 22788 216588 22840
rect 216640 22828 216646 22840
rect 246298 22828 246304 22840
rect 216640 22800 246304 22828
rect 216640 22788 216646 22800
rect 246298 22788 246304 22800
rect 246356 22788 246362 22840
rect 32398 22720 32404 22772
rect 32456 22760 32462 22772
rect 178126 22760 178132 22772
rect 32456 22732 178132 22760
rect 32456 22720 32462 22732
rect 178126 22720 178132 22732
rect 178184 22720 178190 22772
rect 202782 22720 202788 22772
rect 202840 22760 202846 22772
rect 250438 22760 250444 22772
rect 202840 22732 250444 22760
rect 202840 22720 202846 22732
rect 250438 22720 250444 22732
rect 250496 22720 250502 22772
rect 395338 22720 395344 22772
rect 395396 22760 395402 22772
rect 521654 22760 521660 22772
rect 395396 22732 521660 22760
rect 395396 22720 395402 22732
rect 521654 22720 521660 22732
rect 521712 22720 521718 22772
rect 382090 21360 382096 21412
rect 382148 21400 382154 21412
rect 492674 21400 492680 21412
rect 382148 21372 492680 21400
rect 382148 21360 382154 21372
rect 492674 21360 492680 21372
rect 492732 21360 492738 21412
rect 3510 20612 3516 20664
rect 3568 20652 3574 20664
rect 101398 20652 101404 20664
rect 3568 20624 101404 20652
rect 3568 20612 3574 20624
rect 101398 20612 101404 20624
rect 101456 20612 101462 20664
rect 421558 20612 421564 20664
rect 421616 20652 421622 20664
rect 579982 20652 579988 20664
rect 421616 20624 579988 20652
rect 421616 20612 421622 20624
rect 579982 20612 579988 20624
rect 580040 20612 580046 20664
rect 356790 19932 356796 19984
rect 356848 19972 356854 19984
rect 423674 19972 423680 19984
rect 356848 19944 423680 19972
rect 356848 19932 356854 19944
rect 423674 19932 423680 19944
rect 423732 19932 423738 19984
rect 140682 18572 140688 18624
rect 140740 18612 140746 18624
rect 214650 18612 214656 18624
rect 140740 18584 214656 18612
rect 140740 18572 140746 18584
rect 214650 18572 214656 18584
rect 214708 18572 214714 18624
rect 161382 17484 161388 17536
rect 161440 17524 161446 17536
rect 213178 17524 213184 17536
rect 161440 17496 213184 17524
rect 161440 17484 161446 17496
rect 213178 17484 213184 17496
rect 213236 17484 213242 17536
rect 144822 17416 144828 17468
rect 144880 17456 144886 17468
rect 227806 17456 227812 17468
rect 144880 17428 227812 17456
rect 144880 17416 144886 17428
rect 227806 17416 227812 17428
rect 227864 17416 227870 17468
rect 129642 17348 129648 17400
rect 129700 17388 129706 17400
rect 215938 17388 215944 17400
rect 129700 17360 215944 17388
rect 129700 17348 129706 17360
rect 215938 17348 215944 17360
rect 215996 17348 216002 17400
rect 110322 17280 110328 17332
rect 110380 17320 110386 17332
rect 196710 17320 196716 17332
rect 110380 17292 196716 17320
rect 110380 17280 110386 17292
rect 196710 17280 196716 17292
rect 196768 17280 196774 17332
rect 196802 17280 196808 17332
rect 196860 17320 196866 17332
rect 244366 17320 244372 17332
rect 196860 17292 244372 17320
rect 196860 17280 196866 17292
rect 244366 17280 244372 17292
rect 244424 17280 244430 17332
rect 354490 17280 354496 17332
rect 354548 17320 354554 17332
rect 430574 17320 430580 17332
rect 354548 17292 430580 17320
rect 354548 17280 354554 17292
rect 430574 17280 430580 17292
rect 430632 17280 430638 17332
rect 133782 17212 133788 17264
rect 133840 17252 133846 17264
rect 223666 17252 223672 17264
rect 133840 17224 223672 17252
rect 133840 17212 133846 17224
rect 223666 17212 223672 17224
rect 223724 17212 223730 17264
rect 341518 17212 341524 17264
rect 341576 17252 341582 17264
rect 371234 17252 371240 17264
rect 341576 17224 371240 17252
rect 341576 17212 341582 17224
rect 371234 17212 371240 17224
rect 371292 17212 371298 17264
rect 407758 17212 407764 17264
rect 407816 17252 407822 17264
rect 496814 17252 496820 17264
rect 407816 17224 496820 17252
rect 407816 17212 407822 17224
rect 496814 17212 496820 17224
rect 496872 17212 496878 17264
rect 124122 16192 124128 16244
rect 124180 16232 124186 16244
rect 178678 16232 178684 16244
rect 124180 16204 178684 16232
rect 124180 16192 124186 16204
rect 178678 16192 178684 16204
rect 178736 16192 178742 16244
rect 396718 16192 396724 16244
rect 396776 16232 396782 16244
rect 467098 16232 467104 16244
rect 396776 16204 467104 16232
rect 396776 16192 396782 16204
rect 467098 16192 467104 16204
rect 467156 16192 467162 16244
rect 119890 16124 119896 16176
rect 119948 16164 119954 16176
rect 177298 16164 177304 16176
rect 119948 16136 177304 16164
rect 119948 16124 119954 16136
rect 177298 16124 177304 16136
rect 177356 16124 177362 16176
rect 371878 16124 371884 16176
rect 371936 16164 371942 16176
rect 442626 16164 442632 16176
rect 371936 16136 442632 16164
rect 371936 16124 371942 16136
rect 442626 16124 442632 16136
rect 442684 16124 442690 16176
rect 165522 16056 165528 16108
rect 165580 16096 165586 16108
rect 237466 16096 237472 16108
rect 165580 16068 237472 16096
rect 165580 16056 165586 16068
rect 237466 16056 237472 16068
rect 237524 16056 237530 16108
rect 371970 16056 371976 16108
rect 372028 16096 372034 16108
rect 445754 16096 445760 16108
rect 372028 16068 445760 16096
rect 372028 16056 372034 16068
rect 445754 16056 445760 16068
rect 445812 16056 445818 16108
rect 139302 15988 139308 16040
rect 139360 16028 139366 16040
rect 226426 16028 226432 16040
rect 139360 16000 226432 16028
rect 139360 15988 139366 16000
rect 226426 15988 226432 16000
rect 226484 15988 226490 16040
rect 377950 15988 377956 16040
rect 378008 16028 378014 16040
rect 484026 16028 484032 16040
rect 378008 16000 484032 16028
rect 378008 15988 378014 16000
rect 484026 15988 484032 16000
rect 484084 15988 484090 16040
rect 92382 15920 92388 15972
rect 92440 15960 92446 15972
rect 204898 15960 204904 15972
rect 92440 15932 204904 15960
rect 92440 15920 92446 15932
rect 204898 15920 204904 15932
rect 204956 15920 204962 15972
rect 417418 15920 417424 15972
rect 417476 15960 417482 15972
rect 525426 15960 525432 15972
rect 417476 15932 525432 15960
rect 417476 15920 417482 15932
rect 525426 15920 525432 15932
rect 525484 15920 525490 15972
rect 45462 15852 45468 15904
rect 45520 15892 45526 15904
rect 181438 15892 181444 15904
rect 45520 15864 181444 15892
rect 45520 15852 45526 15864
rect 181438 15852 181444 15864
rect 181496 15852 181502 15904
rect 205082 15852 205088 15904
rect 205140 15892 205146 15904
rect 248690 15892 248696 15904
rect 205140 15864 248696 15892
rect 205140 15852 205146 15864
rect 248690 15852 248696 15864
rect 248748 15852 248754 15904
rect 388990 15852 388996 15904
rect 389048 15892 389054 15904
rect 508866 15892 508872 15904
rect 389048 15864 508872 15892
rect 389048 15852 389054 15864
rect 508866 15852 508872 15864
rect 508924 15852 508930 15904
rect 357342 14764 357348 14816
rect 357400 14804 357406 14816
rect 437474 14804 437480 14816
rect 357400 14776 437480 14804
rect 357400 14764 357406 14776
rect 437474 14764 437480 14776
rect 437532 14764 437538 14816
rect 117222 14696 117228 14748
rect 117280 14736 117286 14748
rect 184382 14736 184388 14748
rect 117280 14708 184388 14736
rect 117280 14696 117286 14708
rect 184382 14696 184388 14708
rect 184440 14696 184446 14748
rect 406470 14696 406476 14748
rect 406528 14736 406534 14748
rect 490006 14736 490012 14748
rect 406528 14708 490012 14736
rect 406528 14696 406534 14708
rect 490006 14696 490012 14708
rect 490064 14696 490070 14748
rect 166902 14628 166908 14680
rect 166960 14668 166966 14680
rect 237374 14668 237380 14680
rect 166960 14640 237380 14668
rect 166960 14628 166966 14640
rect 237374 14628 237380 14640
rect 237432 14628 237438 14680
rect 318150 14628 318156 14680
rect 318208 14668 318214 14680
rect 341978 14668 341984 14680
rect 318208 14640 341984 14668
rect 318208 14628 318214 14640
rect 341978 14628 341984 14640
rect 342036 14628 342042 14680
rect 418890 14628 418896 14680
rect 418948 14668 418954 14680
rect 511258 14668 511264 14680
rect 418948 14640 511264 14668
rect 418948 14628 418954 14640
rect 511258 14628 511264 14640
rect 511316 14628 511322 14680
rect 126882 14560 126888 14612
rect 126940 14600 126946 14612
rect 219710 14600 219716 14612
rect 126940 14572 219716 14600
rect 126940 14560 126946 14572
rect 219710 14560 219716 14572
rect 219768 14560 219774 14612
rect 324130 14560 324136 14612
rect 324188 14600 324194 14612
rect 358262 14600 358268 14612
rect 324188 14572 358268 14600
rect 324188 14560 324194 14572
rect 358262 14560 358268 14572
rect 358320 14560 358326 14612
rect 390370 14560 390376 14612
rect 390428 14600 390434 14612
rect 513558 14600 513564 14612
rect 390428 14572 513564 14600
rect 390428 14560 390434 14572
rect 513558 14560 513564 14572
rect 513616 14560 513622 14612
rect 85482 14492 85488 14544
rect 85540 14532 85546 14544
rect 201770 14532 201776 14544
rect 85540 14504 201776 14532
rect 85540 14492 85546 14504
rect 201770 14492 201776 14504
rect 201828 14492 201834 14544
rect 238018 14492 238024 14544
rect 238076 14532 238082 14544
rect 263686 14532 263692 14544
rect 238076 14504 263692 14532
rect 238076 14492 238082 14504
rect 263686 14492 263692 14504
rect 263744 14492 263750 14544
rect 321278 14492 321284 14544
rect 321336 14532 321342 14544
rect 356330 14532 356336 14544
rect 321336 14504 356336 14532
rect 321336 14492 321342 14504
rect 356330 14492 356336 14504
rect 356388 14492 356394 14544
rect 361022 14492 361028 14544
rect 361080 14532 361086 14544
rect 377674 14532 377680 14544
rect 361080 14504 377680 14532
rect 361080 14492 361086 14504
rect 377674 14492 377680 14504
rect 377732 14492 377738 14544
rect 395890 14492 395896 14544
rect 395948 14532 395954 14544
rect 522298 14532 522304 14544
rect 395948 14504 522304 14532
rect 395948 14492 395954 14504
rect 522298 14492 522304 14504
rect 522356 14492 522362 14544
rect 19242 14424 19248 14476
rect 19300 14464 19306 14476
rect 172698 14464 172704 14476
rect 19300 14436 172704 14464
rect 19300 14424 19306 14436
rect 172698 14424 172704 14436
rect 172756 14424 172762 14476
rect 202138 14424 202144 14476
rect 202196 14464 202202 14476
rect 245746 14464 245752 14476
rect 202196 14436 245752 14464
rect 202196 14424 202202 14436
rect 245746 14424 245752 14436
rect 245804 14424 245810 14476
rect 246942 14424 246948 14476
rect 247000 14464 247006 14476
rect 273346 14464 273352 14476
rect 247000 14436 273352 14464
rect 247000 14424 247006 14436
rect 273346 14424 273352 14436
rect 273404 14424 273410 14476
rect 329650 14424 329656 14476
rect 329708 14464 329714 14476
rect 367922 14464 367928 14476
rect 329708 14436 367928 14464
rect 329708 14424 329714 14436
rect 367922 14424 367928 14436
rect 367980 14424 367986 14476
rect 393130 14424 393136 14476
rect 393188 14464 393194 14476
rect 520274 14464 520280 14476
rect 393188 14436 520280 14464
rect 393188 14424 393194 14436
rect 520274 14424 520280 14436
rect 520332 14424 520338 14476
rect 145926 13132 145932 13184
rect 145984 13172 145990 13184
rect 229186 13172 229192 13184
rect 145984 13144 229192 13172
rect 145984 13132 145990 13144
rect 229186 13132 229192 13144
rect 229244 13132 229250 13184
rect 131022 13064 131028 13116
rect 131080 13104 131086 13116
rect 222286 13104 222292 13116
rect 131080 13076 222292 13104
rect 131080 13064 131086 13076
rect 222286 13064 222292 13076
rect 222344 13064 222350 13116
rect 251082 13064 251088 13116
rect 251140 13104 251146 13116
rect 274818 13104 274824 13116
rect 251140 13076 274824 13104
rect 251140 13064 251146 13076
rect 274818 13064 274824 13076
rect 274876 13064 274882 13116
rect 358722 13064 358728 13116
rect 358780 13104 358786 13116
rect 441522 13104 441528 13116
rect 358780 13076 441528 13104
rect 358780 13064 358786 13076
rect 441522 13064 441528 13076
rect 441580 13064 441586 13116
rect 325418 11840 325424 11892
rect 325476 11840 325482 11892
rect 325436 11812 325464 11840
rect 363506 11812 363512 11824
rect 325436 11784 363512 11812
rect 363506 11772 363512 11784
rect 363564 11772 363570 11824
rect 379330 11772 379336 11824
rect 379388 11812 379394 11824
rect 487154 11812 487160 11824
rect 379388 11784 487160 11812
rect 379388 11772 379394 11784
rect 487154 11772 487160 11784
rect 487212 11772 487218 11824
rect 328362 11704 328368 11756
rect 328420 11744 328426 11756
rect 370130 11744 370136 11756
rect 328420 11716 370136 11744
rect 328420 11704 328426 11716
rect 370130 11704 370136 11716
rect 370188 11704 370194 11756
rect 382182 11704 382188 11756
rect 382240 11744 382246 11756
rect 494698 11744 494704 11756
rect 382240 11716 494704 11744
rect 382240 11704 382246 11716
rect 494698 11704 494704 11716
rect 494756 11704 494762 11756
rect 358170 10412 358176 10464
rect 358228 10452 358234 10464
rect 433978 10452 433984 10464
rect 358228 10424 433984 10452
rect 358228 10412 358234 10424
rect 433978 10412 433984 10424
rect 434036 10412 434042 10464
rect 367830 10344 367836 10396
rect 367888 10384 367894 10396
rect 403618 10384 403624 10396
rect 367888 10356 403624 10384
rect 367888 10344 367894 10356
rect 403618 10344 403624 10356
rect 403676 10344 403682 10396
rect 403710 10344 403716 10396
rect 403768 10384 403774 10396
rect 482094 10384 482100 10396
rect 403768 10356 482100 10384
rect 403768 10344 403774 10356
rect 482094 10344 482100 10356
rect 482152 10344 482158 10396
rect 363690 10276 363696 10328
rect 363748 10316 363754 10328
rect 375098 10316 375104 10328
rect 363748 10288 375104 10316
rect 363748 10276 363754 10288
rect 375098 10276 375104 10288
rect 375156 10276 375162 10328
rect 473906 10316 473912 10328
rect 383626 10288 473912 10316
rect 374638 10208 374644 10260
rect 374696 10248 374702 10260
rect 383626 10248 383654 10288
rect 473906 10276 473912 10288
rect 473964 10276 473970 10328
rect 374696 10220 383654 10248
rect 374696 10208 374702 10220
rect 175458 9528 175464 9580
rect 175516 9568 175522 9580
rect 241606 9568 241612 9580
rect 175516 9540 241612 9568
rect 175516 9528 175522 9540
rect 241606 9528 241612 9540
rect 241664 9528 241670 9580
rect 171962 9460 171968 9512
rect 172020 9500 172026 9512
rect 240226 9500 240232 9512
rect 172020 9472 240232 9500
rect 172020 9460 172026 9472
rect 240226 9460 240232 9472
rect 240284 9460 240290 9512
rect 136450 9392 136456 9444
rect 136508 9432 136514 9444
rect 214558 9432 214564 9444
rect 136508 9404 214564 9432
rect 136508 9392 136514 9404
rect 214558 9392 214564 9404
rect 214616 9392 214622 9444
rect 135254 9324 135260 9376
rect 135312 9364 135318 9376
rect 223850 9364 223856 9376
rect 135312 9336 223856 9364
rect 135312 9324 135318 9336
rect 223850 9324 223856 9336
rect 223908 9324 223914 9376
rect 350350 9324 350356 9376
rect 350408 9364 350414 9376
rect 420178 9364 420184 9376
rect 350408 9336 420184 9364
rect 350408 9324 350414 9336
rect 420178 9324 420184 9336
rect 420236 9324 420242 9376
rect 131758 9256 131764 9308
rect 131816 9296 131822 9308
rect 222378 9296 222384 9308
rect 131816 9268 222384 9296
rect 131816 9256 131822 9268
rect 222378 9256 222384 9268
rect 222436 9256 222442 9308
rect 353110 9256 353116 9308
rect 353168 9296 353174 9308
rect 427262 9296 427268 9308
rect 353168 9268 427268 9296
rect 353168 9256 353174 9268
rect 427262 9256 427268 9268
rect 427320 9256 427326 9308
rect 77386 9188 77392 9240
rect 77444 9228 77450 9240
rect 198826 9228 198832 9240
rect 77444 9200 198832 9228
rect 77444 9188 77450 9200
rect 198826 9188 198832 9200
rect 198884 9188 198890 9240
rect 385678 9188 385684 9240
rect 385736 9228 385742 9240
rect 460382 9228 460388 9240
rect 385736 9200 460388 9228
rect 385736 9188 385742 9200
rect 460382 9188 460388 9200
rect 460440 9188 460446 9240
rect 73798 9120 73804 9172
rect 73856 9160 73862 9172
rect 197630 9160 197636 9172
rect 73856 9132 197636 9160
rect 73856 9120 73862 9132
rect 197630 9120 197636 9132
rect 197688 9120 197694 9172
rect 360102 9120 360108 9172
rect 360160 9160 360166 9172
rect 445018 9160 445024 9172
rect 360160 9132 445024 9160
rect 360160 9120 360166 9132
rect 445018 9120 445024 9132
rect 445076 9120 445082 9172
rect 70302 9052 70308 9104
rect 70360 9092 70366 9104
rect 196066 9092 196072 9104
rect 70360 9064 196072 9092
rect 70360 9052 70366 9064
rect 196066 9052 196072 9064
rect 196124 9052 196130 9104
rect 377398 9052 377404 9104
rect 377456 9092 377462 9104
rect 478046 9092 478052 9104
rect 377456 9064 478052 9092
rect 377456 9052 377462 9064
rect 478046 9052 478052 9064
rect 478104 9052 478110 9104
rect 66714 8984 66720 9036
rect 66772 9024 66778 9036
rect 194686 9024 194692 9036
rect 66772 8996 194692 9024
rect 66772 8984 66778 8996
rect 194686 8984 194692 8996
rect 194744 8984 194750 9036
rect 376570 8984 376576 9036
rect 376628 9024 376634 9036
rect 480530 9024 480536 9036
rect 376628 8996 480536 9024
rect 376628 8984 376634 8996
rect 480530 8984 480536 8996
rect 480588 8984 480594 9036
rect 482370 8984 482376 9036
rect 482428 9024 482434 9036
rect 518342 9024 518348 9036
rect 482428 8996 518348 9024
rect 482428 8984 482434 8996
rect 518342 8984 518348 8996
rect 518400 8984 518406 9036
rect 63218 8916 63224 8968
rect 63276 8956 63282 8968
rect 193306 8956 193312 8968
rect 63276 8928 193312 8956
rect 63276 8916 63282 8928
rect 193306 8916 193312 8928
rect 193364 8916 193370 8968
rect 383470 8916 383476 8968
rect 383528 8956 383534 8968
rect 498194 8956 498200 8968
rect 383528 8928 498200 8956
rect 383528 8916 383534 8928
rect 498194 8916 498200 8928
rect 498252 8916 498258 8968
rect 108114 8236 108120 8288
rect 108172 8276 108178 8288
rect 212626 8276 212632 8288
rect 108172 8248 212632 8276
rect 108172 8236 108178 8248
rect 212626 8236 212632 8248
rect 212684 8236 212690 8288
rect 401318 8236 401324 8288
rect 401376 8276 401382 8288
rect 538398 8276 538404 8288
rect 401376 8248 538404 8276
rect 401376 8236 401382 8248
rect 538398 8236 538404 8248
rect 538456 8236 538462 8288
rect 104526 8168 104532 8220
rect 104584 8208 104590 8220
rect 211338 8208 211344 8220
rect 104584 8180 211344 8208
rect 104584 8168 104590 8180
rect 211338 8168 211344 8180
rect 211396 8168 211402 8220
rect 402790 8168 402796 8220
rect 402848 8208 402854 8220
rect 541986 8208 541992 8220
rect 402848 8180 541992 8208
rect 402848 8168 402854 8180
rect 541986 8168 541992 8180
rect 542044 8168 542050 8220
rect 101030 8100 101036 8152
rect 101088 8140 101094 8152
rect 209958 8140 209964 8152
rect 101088 8112 209964 8140
rect 101088 8100 101094 8112
rect 209958 8100 209964 8112
rect 210016 8100 210022 8152
rect 404170 8100 404176 8152
rect 404228 8140 404234 8152
rect 545482 8140 545488 8152
rect 404228 8112 545488 8140
rect 404228 8100 404234 8112
rect 545482 8100 545488 8112
rect 545540 8100 545546 8152
rect 97442 8032 97448 8084
rect 97500 8072 97506 8084
rect 207198 8072 207204 8084
rect 97500 8044 207204 8072
rect 97500 8032 97506 8044
rect 207198 8032 207204 8044
rect 207256 8032 207262 8084
rect 405550 8032 405556 8084
rect 405608 8072 405614 8084
rect 549070 8072 549076 8084
rect 405608 8044 549076 8072
rect 405608 8032 405614 8044
rect 549070 8032 549076 8044
rect 549128 8032 549134 8084
rect 93946 7964 93952 8016
rect 94004 8004 94010 8016
rect 205818 8004 205824 8016
rect 94004 7976 205824 8004
rect 94004 7964 94010 7976
rect 205818 7964 205824 7976
rect 205876 7964 205882 8016
rect 408310 7964 408316 8016
rect 408368 8004 408374 8016
rect 552658 8004 552664 8016
rect 408368 7976 552664 8004
rect 408368 7964 408374 7976
rect 552658 7964 552664 7976
rect 552716 7964 552722 8016
rect 90358 7896 90364 7948
rect 90416 7936 90422 7948
rect 204346 7936 204352 7948
rect 90416 7908 204352 7936
rect 90416 7896 90422 7908
rect 204346 7896 204352 7908
rect 204404 7896 204410 7948
rect 409690 7896 409696 7948
rect 409748 7936 409754 7948
rect 556154 7936 556160 7948
rect 409748 7908 556160 7936
rect 409748 7896 409754 7908
rect 556154 7896 556160 7908
rect 556212 7896 556218 7948
rect 86862 7828 86868 7880
rect 86920 7868 86926 7880
rect 203058 7868 203064 7880
rect 86920 7840 203064 7868
rect 86920 7828 86926 7840
rect 203058 7828 203064 7840
rect 203116 7828 203122 7880
rect 410978 7828 410984 7880
rect 411036 7868 411042 7880
rect 559742 7868 559748 7880
rect 411036 7840 559748 7868
rect 411036 7828 411042 7840
rect 559742 7828 559748 7840
rect 559800 7828 559806 7880
rect 59630 7760 59636 7812
rect 59688 7800 59694 7812
rect 190546 7800 190552 7812
rect 59688 7772 190552 7800
rect 59688 7760 59694 7772
rect 190546 7760 190552 7772
rect 190604 7760 190610 7812
rect 412542 7760 412548 7812
rect 412600 7800 412606 7812
rect 563238 7800 563244 7812
rect 412600 7772 563244 7800
rect 412600 7760 412606 7772
rect 563238 7760 563244 7772
rect 563296 7760 563302 7812
rect 56042 7692 56048 7744
rect 56100 7732 56106 7744
rect 189350 7732 189356 7744
rect 56100 7704 189356 7732
rect 56100 7692 56106 7704
rect 189350 7692 189356 7704
rect 189408 7692 189414 7744
rect 413738 7692 413744 7744
rect 413796 7732 413802 7744
rect 566826 7732 566832 7744
rect 413796 7704 566832 7732
rect 413796 7692 413802 7704
rect 566826 7692 566832 7704
rect 566884 7692 566890 7744
rect 52546 7624 52552 7676
rect 52604 7664 52610 7676
rect 187786 7664 187792 7676
rect 52604 7636 187792 7664
rect 52604 7624 52610 7636
rect 187786 7624 187792 7636
rect 187844 7624 187850 7676
rect 415210 7624 415216 7676
rect 415268 7664 415274 7676
rect 570322 7664 570328 7676
rect 415268 7636 570328 7664
rect 415268 7624 415274 7636
rect 570322 7624 570328 7636
rect 570380 7624 570386 7676
rect 48958 7556 48964 7608
rect 49016 7596 49022 7608
rect 186406 7596 186412 7608
rect 49016 7568 186412 7596
rect 49016 7556 49022 7568
rect 186406 7556 186412 7568
rect 186464 7556 186470 7608
rect 416590 7556 416596 7608
rect 416648 7596 416654 7608
rect 573910 7596 573916 7608
rect 416648 7568 573916 7596
rect 416648 7556 416654 7568
rect 573910 7556 573916 7568
rect 573968 7556 573974 7608
rect 111610 7488 111616 7540
rect 111668 7528 111674 7540
rect 214098 7528 214104 7540
rect 111668 7500 214104 7528
rect 111668 7488 111674 7500
rect 214098 7488 214104 7500
rect 214156 7488 214162 7540
rect 400030 7488 400036 7540
rect 400088 7528 400094 7540
rect 534902 7528 534908 7540
rect 400088 7500 534908 7528
rect 400088 7488 400094 7500
rect 534902 7488 534908 7500
rect 534960 7488 534966 7540
rect 115198 7420 115204 7472
rect 115256 7460 115262 7472
rect 215570 7460 215576 7472
rect 115256 7432 215576 7460
rect 115256 7420 115262 7432
rect 215570 7420 215576 7432
rect 215628 7420 215634 7472
rect 398742 7420 398748 7472
rect 398800 7460 398806 7472
rect 531314 7460 531320 7472
rect 398800 7432 531320 7460
rect 398800 7420 398806 7432
rect 531314 7420 531320 7432
rect 531372 7420 531378 7472
rect 118786 7352 118792 7404
rect 118844 7392 118850 7404
rect 216766 7392 216772 7404
rect 118844 7364 216772 7392
rect 118844 7352 118850 7364
rect 216766 7352 216772 7364
rect 216824 7352 216830 7404
rect 397270 7352 397276 7404
rect 397328 7392 397334 7404
rect 527818 7392 527824 7404
rect 397328 7364 527824 7392
rect 397328 7352 397334 7364
rect 527818 7352 527824 7364
rect 527876 7352 527882 7404
rect 122282 7284 122288 7336
rect 122340 7324 122346 7336
rect 218238 7324 218244 7336
rect 122340 7296 218244 7324
rect 122340 7284 122346 7296
rect 218238 7284 218244 7296
rect 218296 7284 218302 7336
rect 355962 7284 355968 7336
rect 356020 7324 356026 7336
rect 435542 7324 435548 7336
rect 356020 7296 435548 7324
rect 356020 7284 356026 7296
rect 435542 7284 435548 7296
rect 435600 7284 435606 7336
rect 149514 7216 149520 7268
rect 149572 7256 149578 7268
rect 230658 7256 230664 7268
rect 149572 7228 230664 7256
rect 149572 7216 149578 7228
rect 230658 7216 230664 7228
rect 230716 7216 230722 7268
rect 354582 7216 354588 7268
rect 354640 7256 354646 7268
rect 432046 7256 432052 7268
rect 354640 7228 432052 7256
rect 354640 7216 354646 7228
rect 432046 7216 432052 7228
rect 432104 7216 432110 7268
rect 153010 7148 153016 7200
rect 153068 7188 153074 7200
rect 232130 7188 232136 7200
rect 153068 7160 232136 7188
rect 153068 7148 153074 7160
rect 232130 7148 232136 7160
rect 232188 7148 232194 7200
rect 353202 7148 353208 7200
rect 353260 7188 353266 7200
rect 428458 7188 428464 7200
rect 353260 7160 428464 7188
rect 353260 7148 353266 7160
rect 428458 7148 428464 7160
rect 428516 7148 428522 7200
rect 156598 7080 156604 7132
rect 156656 7120 156662 7132
rect 233326 7120 233332 7132
rect 156656 7092 233332 7120
rect 156656 7080 156662 7092
rect 233326 7080 233332 7092
rect 233384 7080 233390 7132
rect 351822 7080 351828 7132
rect 351880 7120 351886 7132
rect 424962 7120 424968 7132
rect 351880 7092 424968 7120
rect 351880 7080 351886 7092
rect 424962 7080 424968 7092
rect 425020 7080 425026 7132
rect 160094 7012 160100 7064
rect 160152 7052 160158 7064
rect 234798 7052 234804 7064
rect 160152 7024 234804 7052
rect 160152 7012 160158 7024
rect 234798 7012 234804 7024
rect 234856 7012 234862 7064
rect 350442 7012 350448 7064
rect 350500 7052 350506 7064
rect 421374 7052 421380 7064
rect 350500 7024 421380 7052
rect 350500 7012 350506 7024
rect 421374 7012 421380 7024
rect 421432 7012 421438 7064
rect 83274 6808 83280 6860
rect 83332 6848 83338 6860
rect 201678 6848 201684 6860
rect 83332 6820 201684 6848
rect 83332 6808 83338 6820
rect 201678 6808 201684 6820
rect 201736 6808 201742 6860
rect 447778 6808 447784 6860
rect 447836 6848 447842 6860
rect 580166 6848 580172 6860
rect 447836 6820 580172 6848
rect 447836 6808 447842 6820
rect 580166 6808 580172 6820
rect 580224 6808 580230 6860
rect 79686 6740 79692 6792
rect 79744 6780 79750 6792
rect 200114 6780 200120 6792
rect 79744 6752 200120 6780
rect 79744 6740 79750 6752
rect 200114 6740 200120 6752
rect 200172 6740 200178 6792
rect 376662 6740 376668 6792
rect 376720 6780 376726 6792
rect 481726 6780 481732 6792
rect 376720 6752 481732 6780
rect 376720 6740 376726 6752
rect 481726 6740 481732 6752
rect 481784 6740 481790 6792
rect 44266 6672 44272 6724
rect 44324 6712 44330 6724
rect 185026 6712 185032 6724
rect 44324 6684 185032 6712
rect 44324 6672 44330 6684
rect 185026 6672 185032 6684
rect 185084 6672 185090 6724
rect 378042 6672 378048 6724
rect 378100 6712 378106 6724
rect 485222 6712 485228 6724
rect 378100 6684 485228 6712
rect 378100 6672 378106 6684
rect 485222 6672 485228 6684
rect 485280 6672 485286 6724
rect 40678 6604 40684 6656
rect 40736 6644 40742 6656
rect 182266 6644 182272 6656
rect 40736 6616 182272 6644
rect 40736 6604 40742 6616
rect 182266 6604 182272 6616
rect 182324 6604 182330 6656
rect 205174 6604 205180 6656
rect 205232 6644 205238 6656
rect 254026 6644 254032 6656
rect 205232 6616 254032 6644
rect 205232 6604 205238 6616
rect 254026 6604 254032 6616
rect 254084 6604 254090 6656
rect 379422 6604 379428 6656
rect 379480 6644 379486 6656
rect 488810 6644 488816 6656
rect 379480 6616 488816 6644
rect 379480 6604 379486 6616
rect 488810 6604 488816 6616
rect 488868 6604 488874 6656
rect 37182 6536 37188 6588
rect 37240 6576 37246 6588
rect 180978 6576 180984 6588
rect 37240 6548 180984 6576
rect 37240 6536 37246 6548
rect 180978 6536 180984 6548
rect 181036 6536 181042 6588
rect 201494 6536 201500 6588
rect 201552 6576 201558 6588
rect 252830 6576 252836 6588
rect 201552 6548 252836 6576
rect 201552 6536 201558 6548
rect 252830 6536 252836 6548
rect 252888 6536 252894 6588
rect 380710 6536 380716 6588
rect 380768 6576 380774 6588
rect 492306 6576 492312 6588
rect 380768 6548 492312 6576
rect 380768 6536 380774 6548
rect 492306 6536 492312 6548
rect 492364 6536 492370 6588
rect 33594 6468 33600 6520
rect 33652 6508 33658 6520
rect 179506 6508 179512 6520
rect 33652 6480 179512 6508
rect 33652 6468 33658 6480
rect 179506 6468 179512 6480
rect 179564 6468 179570 6520
rect 197906 6468 197912 6520
rect 197964 6508 197970 6520
rect 251266 6508 251272 6520
rect 197964 6480 251272 6508
rect 197964 6468 197970 6480
rect 251266 6468 251272 6480
rect 251324 6468 251330 6520
rect 383562 6468 383568 6520
rect 383620 6508 383626 6520
rect 495894 6508 495900 6520
rect 383620 6480 495900 6508
rect 383620 6468 383626 6480
rect 495894 6468 495900 6480
rect 495952 6468 495958 6520
rect 30098 6400 30104 6452
rect 30156 6440 30162 6452
rect 178218 6440 178224 6452
rect 30156 6412 178224 6440
rect 30156 6400 30162 6412
rect 178218 6400 178224 6412
rect 178276 6400 178282 6452
rect 194410 6400 194416 6452
rect 194468 6440 194474 6452
rect 249886 6440 249892 6452
rect 194468 6412 249892 6440
rect 194468 6400 194474 6412
rect 249886 6400 249892 6412
rect 249944 6400 249950 6452
rect 384942 6400 384948 6452
rect 385000 6440 385006 6452
rect 499390 6440 499396 6452
rect 385000 6412 499396 6440
rect 385000 6400 385006 6412
rect 499390 6400 499396 6412
rect 499448 6400 499454 6452
rect 26510 6332 26516 6384
rect 26568 6372 26574 6384
rect 176930 6372 176936 6384
rect 26568 6344 176936 6372
rect 26568 6332 26574 6344
rect 176930 6332 176936 6344
rect 176988 6332 176994 6384
rect 190822 6332 190828 6384
rect 190880 6372 190886 6384
rect 248506 6372 248512 6384
rect 190880 6344 248512 6372
rect 190880 6332 190886 6344
rect 248506 6332 248512 6344
rect 248564 6332 248570 6384
rect 386322 6332 386328 6384
rect 386380 6372 386386 6384
rect 502978 6372 502984 6384
rect 386380 6344 502984 6372
rect 386380 6332 386386 6344
rect 502978 6332 502984 6344
rect 503036 6332 503042 6384
rect 21818 6264 21824 6316
rect 21876 6304 21882 6316
rect 175366 6304 175372 6316
rect 21876 6276 175372 6304
rect 21876 6264 21882 6276
rect 175366 6264 175372 6276
rect 175424 6264 175430 6316
rect 187326 6264 187332 6316
rect 187384 6304 187390 6316
rect 247218 6304 247224 6316
rect 187384 6276 247224 6304
rect 187384 6264 187390 6276
rect 247218 6264 247224 6276
rect 247276 6264 247282 6316
rect 338758 6264 338764 6316
rect 338816 6304 338822 6316
rect 352834 6304 352840 6316
rect 338816 6276 352840 6304
rect 338816 6264 338822 6276
rect 352834 6264 352840 6276
rect 352892 6264 352898 6316
rect 387610 6264 387616 6316
rect 387668 6304 387674 6316
rect 506474 6304 506480 6316
rect 387668 6276 506480 6304
rect 387668 6264 387674 6276
rect 506474 6264 506480 6276
rect 506532 6264 506538 6316
rect 8754 6196 8760 6248
rect 8812 6236 8818 6248
rect 168374 6236 168380 6248
rect 8812 6208 168380 6236
rect 8812 6196 8818 6208
rect 168374 6196 168380 6208
rect 168432 6196 168438 6248
rect 170766 6196 170772 6248
rect 170824 6236 170830 6248
rect 240318 6236 240324 6248
rect 170824 6208 240324 6236
rect 170824 6196 170830 6208
rect 240318 6196 240324 6208
rect 240376 6196 240382 6248
rect 340138 6196 340144 6248
rect 340196 6236 340202 6248
rect 366910 6236 366916 6248
rect 340196 6208 366916 6236
rect 340196 6196 340202 6208
rect 366910 6196 366916 6208
rect 366968 6196 366974 6248
rect 389082 6196 389088 6248
rect 389140 6236 389146 6248
rect 510062 6236 510068 6248
rect 389140 6208 510068 6236
rect 389140 6196 389146 6208
rect 510062 6196 510068 6208
rect 510120 6196 510126 6248
rect 4062 6128 4068 6180
rect 4120 6168 4126 6180
rect 167086 6168 167092 6180
rect 4120 6140 167092 6168
rect 4120 6128 4126 6140
rect 167086 6128 167092 6140
rect 167144 6128 167150 6180
rect 167178 6128 167184 6180
rect 167236 6168 167242 6180
rect 238754 6168 238760 6180
rect 167236 6140 238760 6168
rect 167236 6128 167242 6140
rect 238754 6128 238760 6140
rect 238812 6128 238818 6180
rect 317230 6128 317236 6180
rect 317288 6168 317294 6180
rect 345750 6168 345756 6180
rect 317288 6140 345756 6168
rect 317288 6128 317294 6140
rect 345750 6128 345756 6140
rect 345808 6128 345814 6180
rect 367738 6128 367744 6180
rect 367796 6168 367802 6180
rect 396534 6168 396540 6180
rect 367796 6140 396540 6168
rect 367796 6128 367802 6140
rect 396534 6128 396540 6140
rect 396592 6128 396598 6180
rect 417970 6128 417976 6180
rect 418028 6168 418034 6180
rect 577406 6168 577412 6180
rect 418028 6140 577412 6168
rect 418028 6128 418034 6140
rect 577406 6128 577412 6140
rect 577464 6128 577470 6180
rect 128170 6060 128176 6112
rect 128228 6100 128234 6112
rect 220906 6100 220912 6112
rect 128228 6072 220912 6100
rect 128228 6060 128234 6072
rect 220906 6060 220912 6072
rect 220964 6060 220970 6112
rect 372522 6060 372528 6112
rect 372580 6100 372586 6112
rect 473446 6100 473452 6112
rect 372580 6072 473452 6100
rect 372580 6060 372586 6072
rect 473446 6060 473452 6072
rect 473504 6060 473510 6112
rect 141234 5992 141240 6044
rect 141292 6032 141298 6044
rect 226518 6032 226524 6044
rect 141292 6004 226524 6032
rect 141292 5992 141298 6004
rect 226518 5992 226524 6004
rect 226576 5992 226582 6044
rect 375190 5992 375196 6044
rect 375248 6032 375254 6044
rect 476942 6032 476948 6044
rect 375248 6004 476948 6032
rect 375248 5992 375254 6004
rect 476942 5992 476948 6004
rect 477000 5992 477006 6044
rect 144730 5924 144736 5976
rect 144788 5964 144794 5976
rect 227990 5964 227996 5976
rect 144788 5936 227996 5964
rect 144788 5924 144794 5936
rect 227990 5924 227996 5936
rect 228048 5924 228054 5976
rect 371142 5924 371148 5976
rect 371200 5964 371206 5976
rect 469858 5964 469864 5976
rect 371200 5936 469864 5964
rect 371200 5924 371206 5936
rect 469858 5924 469864 5936
rect 469916 5924 469922 5976
rect 148318 5856 148324 5908
rect 148376 5896 148382 5908
rect 230566 5896 230572 5908
rect 148376 5868 230572 5896
rect 148376 5856 148382 5868
rect 230566 5856 230572 5868
rect 230624 5856 230630 5908
rect 369762 5856 369768 5908
rect 369820 5896 369826 5908
rect 466270 5896 466276 5908
rect 369820 5868 466276 5896
rect 369820 5856 369826 5868
rect 466270 5856 466276 5868
rect 466328 5856 466334 5908
rect 151814 5788 151820 5840
rect 151872 5828 151878 5840
rect 231946 5828 231952 5840
rect 151872 5800 231952 5828
rect 151872 5788 151878 5800
rect 231946 5788 231952 5800
rect 232004 5788 232010 5840
rect 368382 5788 368388 5840
rect 368440 5828 368446 5840
rect 462774 5828 462780 5840
rect 368440 5800 462780 5828
rect 368440 5788 368446 5800
rect 462774 5788 462780 5800
rect 462832 5788 462838 5840
rect 155402 5720 155408 5772
rect 155460 5760 155466 5772
rect 233234 5760 233240 5772
rect 155460 5732 233240 5760
rect 155460 5720 155466 5732
rect 233234 5720 233240 5732
rect 233292 5720 233298 5772
rect 367002 5720 367008 5772
rect 367060 5760 367066 5772
rect 459186 5760 459192 5772
rect 367060 5732 459192 5760
rect 367060 5720 367066 5732
rect 459186 5720 459192 5732
rect 459244 5720 459250 5772
rect 158898 5652 158904 5704
rect 158956 5692 158962 5704
rect 234706 5692 234712 5704
rect 158956 5664 234712 5692
rect 158956 5652 158962 5664
rect 234706 5652 234712 5664
rect 234764 5652 234770 5704
rect 365622 5652 365628 5704
rect 365680 5692 365686 5704
rect 455690 5692 455696 5704
rect 365680 5664 455696 5692
rect 365680 5652 365686 5664
rect 455690 5652 455696 5664
rect 455748 5652 455754 5704
rect 163682 5584 163688 5636
rect 163740 5624 163746 5636
rect 236270 5624 236276 5636
rect 163740 5596 236276 5624
rect 163740 5584 163746 5596
rect 236270 5584 236276 5596
rect 236328 5584 236334 5636
rect 364242 5584 364248 5636
rect 364300 5624 364306 5636
rect 452102 5624 452108 5636
rect 364300 5596 452108 5624
rect 364300 5584 364306 5596
rect 452102 5584 452108 5596
rect 452160 5584 452166 5636
rect 62022 5448 62028 5500
rect 62080 5488 62086 5500
rect 191926 5488 191932 5500
rect 62080 5460 191932 5488
rect 62080 5448 62086 5460
rect 191926 5448 191932 5460
rect 191984 5448 191990 5500
rect 221550 5448 221556 5500
rect 221608 5488 221614 5500
rect 262398 5488 262404 5500
rect 221608 5460 262404 5488
rect 221608 5448 221614 5460
rect 262398 5448 262404 5460
rect 262456 5448 262462 5500
rect 339310 5448 339316 5500
rect 339368 5488 339374 5500
rect 395338 5488 395344 5500
rect 339368 5460 395344 5488
rect 339368 5448 339374 5460
rect 395338 5448 395344 5460
rect 395396 5448 395402 5500
rect 402882 5448 402888 5500
rect 402940 5488 402946 5500
rect 540790 5488 540796 5500
rect 402940 5460 540796 5488
rect 402940 5448 402946 5460
rect 540790 5448 540796 5460
rect 540848 5448 540854 5500
rect 58434 5380 58440 5432
rect 58492 5420 58498 5432
rect 190638 5420 190644 5432
rect 58492 5392 190644 5420
rect 58492 5380 58498 5392
rect 190638 5380 190644 5392
rect 190696 5380 190702 5432
rect 218054 5380 218060 5432
rect 218112 5420 218118 5432
rect 261018 5420 261024 5432
rect 218112 5392 261024 5420
rect 218112 5380 218118 5392
rect 261018 5380 261024 5392
rect 261076 5380 261082 5432
rect 340690 5380 340696 5432
rect 340748 5420 340754 5432
rect 398926 5420 398932 5432
rect 340748 5392 398932 5420
rect 340748 5380 340754 5392
rect 398926 5380 398932 5392
rect 398984 5380 398990 5432
rect 404262 5380 404268 5432
rect 404320 5420 404326 5432
rect 544378 5420 544384 5432
rect 404320 5392 544384 5420
rect 404320 5380 404326 5392
rect 544378 5380 544384 5392
rect 544436 5380 544442 5432
rect 54938 5312 54944 5364
rect 54996 5352 55002 5364
rect 189258 5352 189264 5364
rect 54996 5324 189264 5352
rect 54996 5312 55002 5324
rect 189258 5312 189264 5324
rect 189316 5312 189322 5364
rect 214466 5312 214472 5364
rect 214524 5352 214530 5364
rect 258258 5352 258264 5364
rect 214524 5324 258264 5352
rect 214524 5312 214530 5324
rect 258258 5312 258264 5324
rect 258316 5312 258322 5364
rect 340782 5312 340788 5364
rect 340840 5352 340846 5364
rect 400122 5352 400128 5364
rect 340840 5324 400128 5352
rect 340840 5312 340846 5324
rect 400122 5312 400128 5324
rect 400180 5312 400186 5364
rect 405642 5312 405648 5364
rect 405700 5352 405706 5364
rect 547874 5352 547880 5364
rect 405700 5324 547880 5352
rect 405700 5312 405706 5324
rect 547874 5312 547880 5324
rect 547932 5312 547938 5364
rect 51350 5244 51356 5296
rect 51408 5284 51414 5296
rect 187694 5284 187700 5296
rect 51408 5256 187700 5284
rect 51408 5244 51414 5256
rect 187694 5244 187700 5256
rect 187752 5244 187758 5296
rect 211062 5244 211068 5296
rect 211120 5284 211126 5296
rect 256878 5284 256884 5296
rect 211120 5256 256884 5284
rect 211120 5244 211126 5256
rect 256878 5244 256884 5256
rect 256936 5244 256942 5296
rect 307570 5244 307576 5296
rect 307628 5284 307634 5296
rect 324406 5284 324412 5296
rect 307628 5256 324412 5284
rect 307628 5244 307634 5256
rect 324406 5244 324412 5256
rect 324464 5244 324470 5296
rect 342070 5244 342076 5296
rect 342128 5284 342134 5296
rect 402514 5284 402520 5296
rect 342128 5256 402520 5284
rect 342128 5244 342134 5256
rect 402514 5244 402520 5256
rect 402572 5244 402578 5296
rect 407022 5244 407028 5296
rect 407080 5284 407086 5296
rect 551462 5284 551468 5296
rect 407080 5256 551468 5284
rect 407080 5244 407086 5256
rect 551462 5244 551468 5256
rect 551520 5244 551526 5296
rect 47854 5176 47860 5228
rect 47912 5216 47918 5228
rect 186498 5216 186504 5228
rect 47912 5188 186504 5216
rect 47912 5176 47918 5188
rect 186498 5176 186504 5188
rect 186556 5176 186562 5228
rect 207382 5176 207388 5228
rect 207440 5216 207446 5228
rect 255406 5216 255412 5228
rect 207440 5188 255412 5216
rect 207440 5176 207446 5188
rect 255406 5176 255412 5188
rect 255464 5176 255470 5228
rect 309870 5176 309876 5228
rect 309928 5216 309934 5228
rect 309928 5188 327764 5216
rect 309928 5176 309934 5188
rect 169662 5108 169668 5160
rect 169720 5148 169726 5160
rect 209130 5148 209136 5160
rect 169720 5120 209136 5148
rect 169720 5108 169726 5120
rect 209130 5108 209136 5120
rect 209188 5108 209194 5160
rect 311802 5108 311808 5160
rect 311860 5148 311866 5160
rect 327736 5148 327764 5188
rect 327810 5176 327816 5228
rect 327868 5216 327874 5228
rect 343266 5216 343272 5228
rect 327868 5188 343272 5216
rect 327868 5176 327874 5188
rect 343266 5176 343272 5188
rect 343324 5176 343330 5228
rect 343450 5176 343456 5228
rect 343508 5216 343514 5228
rect 406010 5216 406016 5228
rect 343508 5188 406016 5216
rect 343508 5176 343514 5188
rect 406010 5176 406016 5188
rect 406068 5176 406074 5228
rect 408402 5176 408408 5228
rect 408460 5216 408466 5228
rect 554958 5216 554964 5228
rect 408460 5188 554964 5216
rect 408460 5176 408466 5188
rect 554958 5176 554964 5188
rect 555016 5176 555022 5228
rect 327994 5148 328000 5160
rect 311860 5120 327672 5148
rect 327736 5120 328000 5148
rect 311860 5108 311866 5120
rect 12342 5040 12348 5092
rect 12400 5080 12406 5092
rect 171226 5080 171232 5092
rect 12400 5052 171232 5080
rect 12400 5040 12406 5052
rect 171226 5040 171232 5052
rect 171284 5040 171290 5092
rect 173158 5040 173164 5092
rect 173216 5080 173222 5092
rect 209038 5080 209044 5092
rect 173216 5052 209044 5080
rect 173216 5040 173222 5052
rect 209038 5040 209044 5052
rect 209096 5040 209102 5092
rect 313918 5040 313924 5092
rect 313976 5080 313982 5092
rect 327537 5083 327595 5089
rect 327537 5080 327549 5083
rect 313976 5052 327549 5080
rect 313976 5040 313982 5052
rect 327537 5049 327549 5052
rect 327583 5049 327595 5083
rect 327644 5080 327672 5120
rect 327994 5108 328000 5120
rect 328052 5108 328058 5160
rect 344922 5108 344928 5160
rect 344980 5148 344986 5160
rect 409598 5148 409604 5160
rect 344980 5120 409604 5148
rect 344980 5108 344986 5120
rect 409598 5108 409604 5120
rect 409656 5108 409662 5160
rect 409782 5108 409788 5160
rect 409840 5148 409846 5160
rect 558546 5148 558552 5160
rect 409840 5120 558552 5148
rect 409840 5108 409846 5120
rect 558546 5108 558552 5120
rect 558604 5108 558610 5160
rect 331582 5080 331588 5092
rect 327644 5052 331588 5080
rect 327537 5043 327595 5049
rect 331582 5040 331588 5052
rect 331640 5040 331646 5092
rect 346210 5040 346216 5092
rect 346268 5080 346274 5092
rect 410794 5080 410800 5092
rect 346268 5052 410800 5080
rect 346268 5040 346274 5052
rect 410794 5040 410800 5052
rect 410852 5040 410858 5092
rect 415302 5040 415308 5092
rect 415360 5080 415366 5092
rect 416961 5083 417019 5089
rect 415360 5052 416912 5080
rect 415360 5040 415366 5052
rect 7650 4972 7656 5024
rect 7708 5012 7714 5024
rect 168466 5012 168472 5024
rect 7708 4984 168472 5012
rect 7708 4972 7714 4984
rect 168466 4972 168472 4984
rect 168524 4972 168530 5024
rect 196802 4972 196808 5024
rect 196860 5012 196866 5024
rect 251450 5012 251456 5024
rect 196860 4984 251456 5012
rect 196860 4972 196866 4984
rect 251450 4972 251456 4984
rect 251508 4972 251514 5024
rect 311710 4972 311716 5024
rect 311768 5012 311774 5024
rect 332686 5012 332692 5024
rect 311768 4984 332692 5012
rect 311768 4972 311774 4984
rect 332686 4972 332692 4984
rect 332744 4972 332750 5024
rect 343358 4972 343364 5024
rect 343416 5012 343422 5024
rect 407206 5012 407212 5024
rect 343416 4984 407212 5012
rect 343416 4972 343422 4984
rect 407206 4972 407212 4984
rect 407264 4972 407270 5024
rect 411070 4972 411076 5024
rect 411128 5012 411134 5024
rect 416777 5015 416835 5021
rect 416777 5012 416789 5015
rect 411128 4984 416789 5012
rect 411128 4972 411134 4984
rect 416777 4981 416789 4984
rect 416823 4981 416835 5015
rect 416777 4975 416835 4981
rect 2866 4904 2872 4956
rect 2924 4944 2930 4956
rect 166994 4944 167000 4956
rect 2924 4916 167000 4944
rect 2924 4904 2930 4916
rect 166994 4904 167000 4916
rect 167052 4904 167058 4956
rect 193214 4904 193220 4956
rect 193272 4944 193278 4956
rect 249794 4944 249800 4956
rect 193272 4916 249800 4944
rect 193272 4904 193278 4916
rect 249794 4904 249800 4916
rect 249852 4904 249858 4956
rect 314562 4904 314568 4956
rect 314620 4944 314626 4956
rect 338666 4944 338672 4956
rect 314620 4916 338672 4944
rect 314620 4904 314626 4916
rect 338666 4904 338672 4916
rect 338724 4904 338730 4956
rect 346118 4904 346124 4956
rect 346176 4944 346182 4956
rect 413094 4944 413100 4956
rect 346176 4916 413100 4944
rect 346176 4904 346182 4916
rect 413094 4904 413100 4916
rect 413152 4904 413158 4956
rect 413830 4904 413836 4956
rect 413888 4944 413894 4956
rect 416501 4947 416559 4953
rect 416501 4944 416513 4947
rect 413888 4916 416513 4944
rect 413888 4904 413894 4916
rect 416501 4913 416513 4916
rect 416547 4913 416559 4947
rect 416501 4907 416559 4913
rect 416590 4904 416596 4956
rect 416648 4944 416654 4956
rect 416884 4944 416912 5052
rect 416961 5049 416973 5083
rect 417007 5080 417019 5083
rect 565630 5080 565636 5092
rect 417007 5052 565636 5080
rect 417007 5049 417019 5052
rect 416961 5043 417019 5049
rect 565630 5040 565636 5052
rect 565688 5040 565694 5092
rect 417053 5015 417111 5021
rect 417053 4981 417065 5015
rect 417099 5012 417111 5015
rect 562042 5012 562048 5024
rect 417099 4984 562048 5012
rect 417099 4981 417111 4984
rect 417053 4975 417111 4981
rect 562042 4972 562048 4984
rect 562100 4972 562106 5024
rect 569126 4944 569132 4956
rect 416648 4916 416820 4944
rect 416884 4916 569132 4944
rect 416648 4904 416654 4916
rect 1670 4836 1676 4888
rect 1728 4876 1734 4888
rect 165614 4876 165620 4888
rect 1728 4848 165620 4876
rect 1728 4836 1734 4848
rect 165614 4836 165620 4848
rect 165672 4836 165678 4888
rect 189718 4836 189724 4888
rect 189776 4876 189782 4888
rect 248414 4876 248420 4888
rect 189776 4848 248420 4876
rect 189776 4836 189782 4848
rect 248414 4836 248420 4848
rect 248472 4836 248478 4888
rect 314470 4836 314476 4888
rect 314528 4876 314534 4888
rect 339862 4876 339868 4888
rect 314528 4848 339868 4876
rect 314528 4836 314534 4848
rect 339862 4836 339868 4848
rect 339920 4836 339926 4888
rect 347682 4836 347688 4888
rect 347740 4876 347746 4888
rect 416682 4876 416688 4888
rect 347740 4848 416688 4876
rect 347740 4836 347746 4848
rect 416682 4836 416688 4848
rect 416740 4836 416746 4888
rect 416792 4876 416820 4916
rect 569126 4904 569132 4916
rect 569184 4904 569190 4956
rect 572714 4876 572720 4888
rect 416792 4848 572720 4876
rect 572714 4836 572720 4848
rect 572772 4836 572778 4888
rect 566 4768 572 4820
rect 624 4808 630 4820
rect 165706 4808 165712 4820
rect 624 4780 165712 4808
rect 624 4768 630 4780
rect 165706 4768 165712 4780
rect 165764 4768 165770 4820
rect 174262 4768 174268 4820
rect 174320 4808 174326 4820
rect 241514 4808 241520 4820
rect 174320 4780 241520 4808
rect 174320 4768 174326 4780
rect 241514 4768 241520 4780
rect 241572 4768 241578 4820
rect 318058 4768 318064 4820
rect 318116 4808 318122 4820
rect 346946 4808 346952 4820
rect 318116 4780 346952 4808
rect 318116 4768 318122 4780
rect 346946 4768 346952 4780
rect 347004 4768 347010 4820
rect 349062 4768 349068 4820
rect 349120 4808 349126 4820
rect 417878 4808 417884 4820
rect 349120 4780 417884 4808
rect 349120 4768 349126 4780
rect 417878 4768 417884 4780
rect 417936 4768 417942 4820
rect 418062 4768 418068 4820
rect 418120 4808 418126 4820
rect 576302 4808 576308 4820
rect 418120 4780 576308 4808
rect 418120 4768 418126 4780
rect 576302 4768 576308 4780
rect 576360 4768 576366 4820
rect 65518 4700 65524 4752
rect 65576 4740 65582 4752
rect 193398 4740 193404 4752
rect 65576 4712 193404 4740
rect 65576 4700 65582 4712
rect 193398 4700 193404 4712
rect 193456 4700 193462 4752
rect 200298 4700 200304 4752
rect 200356 4740 200362 4752
rect 252554 4740 252560 4752
rect 200356 4712 252560 4740
rect 200356 4700 200362 4712
rect 252554 4700 252560 4712
rect 252612 4700 252618 4752
rect 327537 4743 327595 4749
rect 327537 4709 327549 4743
rect 327583 4740 327595 4743
rect 334986 4740 334992 4752
rect 327583 4712 334992 4740
rect 327583 4709 327595 4712
rect 327537 4703 327595 4709
rect 334986 4700 334992 4712
rect 335044 4700 335050 4752
rect 337930 4700 337936 4752
rect 337988 4740 337994 4752
rect 393038 4740 393044 4752
rect 337988 4712 393044 4740
rect 337988 4700 337994 4712
rect 393038 4700 393044 4712
rect 393096 4700 393102 4752
rect 401410 4700 401416 4752
rect 401468 4740 401474 4752
rect 537202 4740 537208 4752
rect 401468 4712 537208 4740
rect 401468 4700 401474 4712
rect 537202 4700 537208 4712
rect 537260 4700 537266 4752
rect 72602 4632 72608 4684
rect 72660 4672 72666 4684
rect 197538 4672 197544 4684
rect 72660 4644 197544 4672
rect 72660 4632 72666 4644
rect 197538 4632 197544 4644
rect 197596 4632 197602 4684
rect 203886 4632 203892 4684
rect 203944 4672 203950 4684
rect 254118 4672 254124 4684
rect 203944 4644 254124 4672
rect 203944 4632 203950 4644
rect 254118 4632 254124 4644
rect 254176 4632 254182 4684
rect 335078 4632 335084 4684
rect 335136 4672 335142 4684
rect 388254 4672 388260 4684
rect 335136 4644 388260 4672
rect 335136 4632 335142 4644
rect 388254 4632 388260 4644
rect 388312 4632 388318 4684
rect 400030 4632 400036 4684
rect 400088 4672 400094 4684
rect 533706 4672 533712 4684
rect 400088 4644 533712 4672
rect 400088 4632 400094 4644
rect 533706 4632 533712 4644
rect 533764 4632 533770 4684
rect 69106 4564 69112 4616
rect 69164 4604 69170 4616
rect 194778 4604 194784 4616
rect 69164 4576 194784 4604
rect 69164 4564 69170 4576
rect 194778 4564 194784 4576
rect 194836 4564 194842 4616
rect 338022 4564 338028 4616
rect 338080 4604 338086 4616
rect 391842 4604 391848 4616
rect 338080 4576 391848 4604
rect 338080 4564 338086 4576
rect 391842 4564 391848 4576
rect 391900 4564 391906 4616
rect 397362 4564 397368 4616
rect 397420 4604 397426 4616
rect 530118 4604 530124 4616
rect 397420 4576 530124 4604
rect 397420 4564 397426 4576
rect 530118 4564 530124 4576
rect 530176 4564 530182 4616
rect 76190 4496 76196 4548
rect 76248 4536 76254 4548
rect 198918 4536 198924 4548
rect 76248 4508 198924 4536
rect 76248 4496 76254 4508
rect 198918 4496 198924 4508
rect 198976 4496 198982 4548
rect 335170 4496 335176 4548
rect 335228 4536 335234 4548
rect 385954 4536 385960 4548
rect 335228 4508 385960 4536
rect 335228 4496 335234 4508
rect 385954 4496 385960 4508
rect 386012 4496 386018 4548
rect 395982 4496 395988 4548
rect 396040 4536 396046 4548
rect 526622 4536 526628 4548
rect 396040 4508 526628 4536
rect 396040 4496 396046 4508
rect 526622 4496 526628 4508
rect 526680 4496 526686 4548
rect 126974 4428 126980 4480
rect 127032 4468 127038 4480
rect 220814 4468 220820 4480
rect 127032 4440 220820 4468
rect 127032 4428 127038 4440
rect 220814 4428 220820 4440
rect 220872 4428 220878 4480
rect 333882 4428 333888 4480
rect 333940 4468 333946 4480
rect 384758 4468 384764 4480
rect 333940 4440 384764 4468
rect 333940 4428 333946 4440
rect 384758 4428 384764 4440
rect 384816 4428 384822 4480
rect 394602 4428 394608 4480
rect 394660 4468 394666 4480
rect 523034 4468 523040 4480
rect 394660 4440 523040 4468
rect 394660 4428 394666 4440
rect 523034 4428 523040 4440
rect 523092 4428 523098 4480
rect 150618 4360 150624 4412
rect 150676 4400 150682 4412
rect 230750 4400 230756 4412
rect 150676 4372 230756 4400
rect 150676 4360 150682 4372
rect 230750 4360 230756 4372
rect 230808 4360 230814 4412
rect 332410 4360 332416 4412
rect 332468 4400 332474 4412
rect 381170 4400 381176 4412
rect 332468 4372 381176 4400
rect 332468 4360 332474 4372
rect 381170 4360 381176 4372
rect 381228 4360 381234 4412
rect 393222 4360 393228 4412
rect 393280 4400 393286 4412
rect 519538 4400 519544 4412
rect 393280 4372 519544 4400
rect 393280 4360 393286 4372
rect 519538 4360 519544 4372
rect 519596 4360 519602 4412
rect 154206 4292 154212 4344
rect 154264 4332 154270 4344
rect 231854 4332 231860 4344
rect 154264 4304 231860 4332
rect 154264 4292 154270 4304
rect 231854 4292 231860 4304
rect 231912 4292 231918 4344
rect 332318 4292 332324 4344
rect 332376 4332 332382 4344
rect 378870 4332 378876 4344
rect 332376 4304 378876 4332
rect 332376 4292 332382 4304
rect 378870 4292 378876 4304
rect 378928 4292 378934 4344
rect 391750 4292 391756 4344
rect 391808 4332 391814 4344
rect 515950 4332 515956 4344
rect 391808 4304 515956 4332
rect 391808 4292 391814 4304
rect 515950 4292 515956 4304
rect 516008 4292 516014 4344
rect 157794 4224 157800 4276
rect 157852 4264 157858 4276
rect 234614 4264 234620 4276
rect 157852 4236 234620 4264
rect 157852 4224 157858 4236
rect 234614 4224 234620 4236
rect 234672 4224 234678 4276
rect 367922 4224 367928 4276
rect 367980 4264 367986 4276
rect 367980 4236 369072 4264
rect 367980 4224 367986 4236
rect 17034 4156 17040 4208
rect 17092 4196 17098 4208
rect 172790 4196 172796 4208
rect 17092 4168 172796 4196
rect 17092 4156 17098 4168
rect 172790 4156 172796 4168
rect 172848 4156 172854 4208
rect 177850 4156 177856 4208
rect 177908 4196 177914 4208
rect 224218 4196 224224 4208
rect 177908 4168 224224 4196
rect 177908 4156 177914 4168
rect 224218 4156 224224 4168
rect 224276 4156 224282 4208
rect 347590 4156 347596 4208
rect 347648 4196 347654 4208
rect 368845 4199 368903 4205
rect 368845 4196 368857 4199
rect 347648 4168 368857 4196
rect 347648 4156 347654 4168
rect 368845 4165 368857 4168
rect 368891 4165 368903 4199
rect 368845 4159 368903 4165
rect 61378 4128 61384 4140
rect 26206 4100 61384 4128
rect 11146 4020 11152 4072
rect 11204 4060 11210 4072
rect 18598 4060 18604 4072
rect 11204 4032 18604 4060
rect 11204 4020 11210 4032
rect 18598 4020 18604 4032
rect 18656 4020 18662 4072
rect 20622 4020 20628 4072
rect 20680 4060 20686 4072
rect 26206 4060 26234 4100
rect 61378 4088 61384 4100
rect 61436 4088 61442 4140
rect 64322 4088 64328 4140
rect 64380 4128 64386 4140
rect 184290 4128 184296 4140
rect 64380 4100 184296 4128
rect 64380 4088 64386 4100
rect 184290 4088 184296 4100
rect 184348 4088 184354 4140
rect 242894 4088 242900 4140
rect 242952 4128 242958 4140
rect 267090 4128 267096 4140
rect 242952 4100 267096 4128
rect 242952 4088 242958 4100
rect 267090 4088 267096 4100
rect 267148 4088 267154 4140
rect 281902 4088 281908 4140
rect 281960 4128 281966 4140
rect 288526 4128 288532 4140
rect 281960 4100 288532 4128
rect 281960 4088 281966 4100
rect 288526 4088 288532 4100
rect 288584 4088 288590 4140
rect 296622 4088 296628 4140
rect 296680 4128 296686 4140
rect 297266 4128 297272 4140
rect 296680 4100 297272 4128
rect 296680 4088 296686 4100
rect 297266 4088 297272 4100
rect 297324 4088 297330 4140
rect 303430 4088 303436 4140
rect 303488 4128 303494 4140
rect 312449 4131 312507 4137
rect 312449 4128 312461 4131
rect 303488 4100 312461 4128
rect 303488 4088 303494 4100
rect 312449 4097 312461 4100
rect 312495 4097 312507 4131
rect 312449 4091 312507 4097
rect 312538 4088 312544 4140
rect 312596 4128 312602 4140
rect 316218 4128 316224 4140
rect 312596 4100 316224 4128
rect 312596 4088 312602 4100
rect 316218 4088 316224 4100
rect 316276 4088 316282 4140
rect 331122 4088 331128 4140
rect 331180 4128 331186 4140
rect 368937 4131 368995 4137
rect 368937 4128 368949 4131
rect 331180 4100 368949 4128
rect 331180 4088 331186 4100
rect 368937 4097 368949 4100
rect 368983 4097 368995 4131
rect 369044 4128 369072 4236
rect 390462 4224 390468 4276
rect 390520 4264 390526 4276
rect 512454 4264 512460 4276
rect 390520 4236 512460 4264
rect 390520 4224 390526 4236
rect 512454 4224 512460 4236
rect 512512 4224 512518 4276
rect 369121 4199 369179 4205
rect 369121 4165 369133 4199
rect 369167 4196 369179 4199
rect 414290 4196 414296 4208
rect 369167 4168 414296 4196
rect 369167 4165 369179 4168
rect 369121 4159 369179 4165
rect 414290 4156 414296 4168
rect 414348 4156 414354 4208
rect 490742 4156 490748 4208
rect 490800 4196 490806 4208
rect 490800 4168 491248 4196
rect 490800 4156 490806 4168
rect 374086 4128 374092 4140
rect 369044 4100 374092 4128
rect 368937 4091 368995 4097
rect 374086 4088 374092 4100
rect 374144 4088 374150 4140
rect 381538 4088 381544 4140
rect 381596 4128 381602 4140
rect 472250 4128 472256 4140
rect 381596 4100 472256 4128
rect 381596 4088 381602 4100
rect 472250 4088 472256 4100
rect 472308 4088 472314 4140
rect 489914 4088 489920 4140
rect 489972 4128 489978 4140
rect 491110 4128 491116 4140
rect 489972 4100 491116 4128
rect 489972 4088 489978 4100
rect 491110 4088 491116 4100
rect 491168 4088 491174 4140
rect 491220 4128 491248 4168
rect 582190 4128 582196 4140
rect 491220 4100 582196 4128
rect 582190 4088 582196 4100
rect 582248 4088 582254 4140
rect 20680 4032 26234 4060
rect 20680 4020 20686 4032
rect 35986 4020 35992 4072
rect 36044 4060 36050 4072
rect 51718 4060 51724 4072
rect 36044 4032 51724 4060
rect 36044 4020 36050 4032
rect 51718 4020 51724 4032
rect 51776 4020 51782 4072
rect 53742 4020 53748 4072
rect 53800 4060 53806 4072
rect 57146 4060 57152 4072
rect 53800 4032 57152 4060
rect 53800 4020 53806 4032
rect 57146 4020 57152 4032
rect 57204 4020 57210 4072
rect 57238 4020 57244 4072
rect 57296 4060 57302 4072
rect 184198 4060 184204 4072
rect 57296 4032 184204 4060
rect 57296 4020 57302 4032
rect 184198 4020 184204 4032
rect 184256 4020 184262 4072
rect 228726 4020 228732 4072
rect 228784 4060 228790 4072
rect 242158 4060 242164 4072
rect 228784 4032 242164 4060
rect 228784 4020 228790 4032
rect 242158 4020 242164 4032
rect 242216 4020 242222 4072
rect 244090 4020 244096 4072
rect 244148 4060 244154 4072
rect 258169 4063 258227 4069
rect 244148 4032 258074 4060
rect 244148 4020 244154 4032
rect 50154 3952 50160 4004
rect 50212 3992 50218 4004
rect 176105 3995 176163 4001
rect 50212 3964 176056 3992
rect 50212 3952 50218 3964
rect 46658 3884 46664 3936
rect 46716 3924 46722 3936
rect 175921 3927 175979 3933
rect 175921 3924 175933 3927
rect 46716 3896 175933 3924
rect 46716 3884 46722 3896
rect 175921 3893 175933 3896
rect 175967 3893 175979 3927
rect 175921 3887 175979 3893
rect 39574 3816 39580 3868
rect 39632 3856 39638 3868
rect 176028 3856 176056 3964
rect 176105 3961 176117 3995
rect 176151 3992 176163 3995
rect 185210 3992 185216 4004
rect 176151 3964 185216 3992
rect 176151 3961 176163 3964
rect 176105 3955 176163 3961
rect 185210 3952 185216 3964
rect 185268 3952 185274 4004
rect 232222 3952 232228 4004
rect 232280 3992 232286 4004
rect 253201 3995 253259 4001
rect 253201 3992 253213 3995
rect 232280 3964 253213 3992
rect 232280 3952 232286 3964
rect 253201 3961 253213 3964
rect 253247 3961 253259 3995
rect 258046 3992 258074 4032
rect 258169 4029 258181 4063
rect 258215 4060 258227 4063
rect 266998 4060 267004 4072
rect 258215 4032 267004 4060
rect 258215 4029 258227 4032
rect 258169 4023 258227 4029
rect 266998 4020 267004 4032
rect 267056 4020 267062 4072
rect 306190 4020 306196 4072
rect 306248 4060 306254 4072
rect 319714 4060 319720 4072
rect 306248 4032 319720 4060
rect 306248 4020 306254 4032
rect 319714 4020 319720 4032
rect 319772 4020 319778 4072
rect 329742 4020 329748 4072
rect 329800 4060 329806 4072
rect 372890 4060 372896 4072
rect 329800 4032 372896 4060
rect 329800 4020 329806 4032
rect 372890 4020 372896 4032
rect 372948 4020 372954 4072
rect 375282 4020 375288 4072
rect 375340 4060 375346 4072
rect 479334 4060 479340 4072
rect 375340 4032 479340 4060
rect 375340 4020 375346 4032
rect 479334 4020 479340 4032
rect 479392 4020 479398 4072
rect 486418 4020 486424 4072
rect 486476 4060 486482 4072
rect 578602 4060 578608 4072
rect 486476 4032 578608 4060
rect 486476 4020 486482 4032
rect 578602 4020 578608 4032
rect 578660 4020 578666 4072
rect 269758 3992 269764 4004
rect 258046 3964 269764 3992
rect 253201 3955 253259 3961
rect 269758 3952 269764 3964
rect 269816 3952 269822 4004
rect 306282 3952 306288 4004
rect 306340 3992 306346 4004
rect 320910 3992 320916 4004
rect 306340 3964 320916 3992
rect 306340 3952 306346 3964
rect 320910 3952 320916 3964
rect 320968 3952 320974 4004
rect 332502 3952 332508 4004
rect 332560 3992 332566 4004
rect 379974 3992 379980 4004
rect 332560 3964 379980 3992
rect 332560 3952 332566 3964
rect 379974 3952 379980 3964
rect 380032 3952 380038 4004
rect 399478 3952 399484 4004
rect 399536 3992 399542 4004
rect 532510 3992 532516 4004
rect 399536 3964 532516 3992
rect 399536 3952 399542 3964
rect 532510 3952 532516 3964
rect 532568 3952 532574 4004
rect 192018 3884 192024 3936
rect 192076 3924 192082 3936
rect 205082 3924 205088 3936
rect 192076 3896 205088 3924
rect 192076 3884 192082 3896
rect 205082 3884 205088 3896
rect 205140 3884 205146 3936
rect 225138 3884 225144 3936
rect 225196 3924 225202 3936
rect 238018 3924 238024 3936
rect 225196 3896 238024 3924
rect 225196 3884 225202 3896
rect 238018 3884 238024 3896
rect 238076 3884 238082 3936
rect 241698 3884 241704 3936
rect 241756 3924 241762 3936
rect 269850 3924 269856 3936
rect 241756 3896 269856 3924
rect 241756 3884 241762 3896
rect 269850 3884 269856 3896
rect 269908 3884 269914 3936
rect 300762 3884 300768 3936
rect 300820 3924 300826 3936
rect 306742 3924 306748 3936
rect 300820 3896 306748 3924
rect 300820 3884 300826 3896
rect 306742 3884 306748 3896
rect 306800 3884 306806 3936
rect 312449 3927 312507 3933
rect 312449 3893 312461 3927
rect 312495 3924 312507 3927
rect 313826 3924 313832 3936
rect 312495 3896 313832 3924
rect 312495 3893 312507 3896
rect 312449 3887 312507 3893
rect 313826 3884 313832 3896
rect 313884 3884 313890 3936
rect 325602 3924 325608 3936
rect 313936 3896 325608 3924
rect 182818 3856 182824 3868
rect 39632 3828 175964 3856
rect 176028 3828 182824 3856
rect 39632 3816 39638 3828
rect 19426 3748 19432 3800
rect 19484 3788 19490 3800
rect 29638 3788 29644 3800
rect 19484 3760 29644 3788
rect 19484 3748 19490 3760
rect 29638 3748 29644 3760
rect 29696 3748 29702 3800
rect 32490 3748 32496 3800
rect 32548 3788 32554 3800
rect 175936 3788 175964 3828
rect 182818 3816 182824 3828
rect 182876 3816 182882 3868
rect 199102 3816 199108 3868
rect 199160 3856 199166 3868
rect 206370 3856 206376 3868
rect 199160 3828 206376 3856
rect 199160 3816 199166 3828
rect 206370 3816 206376 3828
rect 206428 3816 206434 3868
rect 219250 3816 219256 3868
rect 219308 3856 219314 3868
rect 232498 3856 232504 3868
rect 219308 3828 232504 3856
rect 219308 3816 219314 3828
rect 232498 3816 232504 3828
rect 232556 3816 232562 3868
rect 237006 3816 237012 3868
rect 237064 3856 237070 3868
rect 258077 3859 258135 3865
rect 258077 3856 258089 3859
rect 237064 3828 258089 3856
rect 237064 3816 237070 3828
rect 258077 3825 258089 3828
rect 258123 3825 258135 3859
rect 264238 3856 264244 3868
rect 258077 3819 258135 3825
rect 258184 3828 264244 3856
rect 182358 3788 182364 3800
rect 32548 3760 175688 3788
rect 175936 3760 182364 3788
rect 32548 3748 32554 3760
rect 67910 3680 67916 3732
rect 67968 3720 67974 3732
rect 76558 3720 76564 3732
rect 67968 3692 76564 3720
rect 67968 3680 67974 3692
rect 76558 3680 76564 3692
rect 76616 3680 76622 3732
rect 80882 3680 80888 3732
rect 80940 3720 80946 3732
rect 81342 3720 81348 3732
rect 80940 3692 81348 3720
rect 80940 3680 80946 3692
rect 81342 3680 81348 3692
rect 81400 3680 81406 3732
rect 84470 3680 84476 3732
rect 84528 3720 84534 3732
rect 85482 3720 85488 3732
rect 84528 3692 85488 3720
rect 84528 3680 84534 3692
rect 85482 3680 85488 3692
rect 85540 3680 85546 3732
rect 91554 3680 91560 3732
rect 91612 3720 91618 3732
rect 92382 3720 92388 3732
rect 91612 3692 92388 3720
rect 91612 3680 91618 3692
rect 92382 3680 92388 3692
rect 92440 3680 92446 3732
rect 92750 3680 92756 3732
rect 92808 3720 92814 3732
rect 94498 3720 94504 3732
rect 92808 3692 94504 3720
rect 92808 3680 92814 3692
rect 94498 3680 94504 3692
rect 94556 3680 94562 3732
rect 98638 3680 98644 3732
rect 98696 3720 98702 3732
rect 99282 3720 99288 3732
rect 98696 3692 99288 3720
rect 98696 3680 98702 3692
rect 99282 3680 99288 3692
rect 99340 3680 99346 3732
rect 99834 3680 99840 3732
rect 99892 3720 99898 3732
rect 101582 3720 101588 3732
rect 99892 3692 101588 3720
rect 99892 3680 99898 3692
rect 101582 3680 101588 3692
rect 101640 3680 101646 3732
rect 102226 3680 102232 3732
rect 102284 3720 102290 3732
rect 103422 3720 103428 3732
rect 102284 3692 103428 3720
rect 102284 3680 102290 3692
rect 103422 3680 103428 3692
rect 103480 3680 103486 3732
rect 105722 3680 105728 3732
rect 105780 3720 105786 3732
rect 106182 3720 106188 3732
rect 105780 3692 106188 3720
rect 105780 3680 105786 3692
rect 106182 3680 106188 3692
rect 106240 3680 106246 3732
rect 106918 3680 106924 3732
rect 106976 3720 106982 3732
rect 107562 3720 107568 3732
rect 106976 3692 107568 3720
rect 106976 3680 106982 3692
rect 107562 3680 107568 3692
rect 107620 3680 107626 3732
rect 109310 3680 109316 3732
rect 109368 3720 109374 3732
rect 110322 3720 110328 3732
rect 109368 3692 110328 3720
rect 109368 3680 109374 3692
rect 110322 3680 110328 3692
rect 110380 3680 110386 3732
rect 114002 3680 114008 3732
rect 114060 3720 114066 3732
rect 114462 3720 114468 3732
rect 114060 3692 114468 3720
rect 114060 3680 114066 3692
rect 114462 3680 114468 3692
rect 114520 3680 114526 3732
rect 116394 3680 116400 3732
rect 116452 3720 116458 3732
rect 117222 3720 117228 3732
rect 116452 3692 117228 3720
rect 116452 3680 116458 3692
rect 117222 3680 117228 3692
rect 117280 3680 117286 3732
rect 123478 3680 123484 3732
rect 123536 3720 123542 3732
rect 124122 3720 124128 3732
rect 123536 3692 124128 3720
rect 123536 3680 123542 3692
rect 124122 3680 124128 3692
rect 124180 3680 124186 3732
rect 124674 3680 124680 3732
rect 124732 3720 124738 3732
rect 125502 3720 125508 3732
rect 124732 3692 125508 3720
rect 124732 3680 124738 3692
rect 125502 3680 125508 3692
rect 125560 3680 125566 3732
rect 125870 3680 125876 3732
rect 125928 3720 125934 3732
rect 126882 3720 126888 3732
rect 125928 3692 126888 3720
rect 125928 3680 125934 3692
rect 126882 3680 126888 3692
rect 126940 3680 126946 3732
rect 130562 3680 130568 3732
rect 130620 3720 130626 3732
rect 131022 3720 131028 3732
rect 130620 3692 131028 3720
rect 130620 3680 130626 3692
rect 131022 3680 131028 3692
rect 131080 3680 131086 3732
rect 132954 3680 132960 3732
rect 133012 3720 133018 3732
rect 133782 3720 133788 3732
rect 133012 3692 133788 3720
rect 133012 3680 133018 3692
rect 133782 3680 133788 3692
rect 133840 3680 133846 3732
rect 134150 3680 134156 3732
rect 134208 3720 134214 3732
rect 135162 3720 135168 3732
rect 134208 3692 135168 3720
rect 134208 3680 134214 3692
rect 135162 3680 135168 3692
rect 135220 3680 135226 3732
rect 138842 3680 138848 3732
rect 138900 3720 138906 3732
rect 139302 3720 139308 3732
rect 138900 3692 139308 3720
rect 138900 3680 138906 3692
rect 139302 3680 139308 3692
rect 139360 3680 139366 3732
rect 140038 3680 140044 3732
rect 140096 3720 140102 3732
rect 140682 3720 140688 3732
rect 140096 3692 140688 3720
rect 140096 3680 140102 3692
rect 140682 3680 140688 3692
rect 140740 3680 140746 3732
rect 142430 3680 142436 3732
rect 142488 3720 142494 3732
rect 143442 3720 143448 3732
rect 142488 3692 143448 3720
rect 142488 3680 142494 3692
rect 143442 3680 143448 3692
rect 143500 3680 143506 3732
rect 143534 3680 143540 3732
rect 143592 3720 143598 3732
rect 144822 3720 144828 3732
rect 143592 3692 144828 3720
rect 143592 3680 143598 3692
rect 144822 3680 144828 3692
rect 144880 3680 144886 3732
rect 147122 3680 147128 3732
rect 147180 3720 147186 3732
rect 147582 3720 147588 3732
rect 147180 3692 147588 3720
rect 147180 3680 147186 3692
rect 147582 3680 147588 3692
rect 147640 3680 147646 3732
rect 164789 3723 164847 3729
rect 164789 3689 164801 3723
rect 164835 3720 164847 3723
rect 168650 3720 168656 3732
rect 164835 3692 168656 3720
rect 164835 3689 164847 3692
rect 164789 3683 164847 3689
rect 168650 3680 168656 3692
rect 168708 3680 168714 3732
rect 24210 3612 24216 3664
rect 24268 3652 24274 3664
rect 175550 3652 175556 3664
rect 24268 3624 175556 3652
rect 24268 3612 24274 3624
rect 175550 3612 175556 3624
rect 175608 3612 175614 3664
rect 175660 3652 175688 3760
rect 182358 3748 182364 3760
rect 182416 3748 182422 3800
rect 184934 3748 184940 3800
rect 184992 3788 184998 3800
rect 202138 3788 202144 3800
rect 184992 3760 202144 3788
rect 184992 3748 184998 3760
rect 202138 3748 202144 3760
rect 202196 3748 202202 3800
rect 223942 3748 223948 3800
rect 224000 3788 224006 3800
rect 256050 3788 256056 3800
rect 224000 3760 256056 3788
rect 224000 3748 224006 3760
rect 256050 3748 256056 3760
rect 256108 3748 256114 3800
rect 258184 3788 258212 3828
rect 264238 3816 264244 3828
rect 264296 3816 264302 3868
rect 300670 3816 300676 3868
rect 300728 3856 300734 3868
rect 307938 3856 307944 3868
rect 300728 3828 307944 3856
rect 300728 3816 300734 3828
rect 307938 3816 307944 3828
rect 307996 3816 308002 3868
rect 309778 3816 309784 3868
rect 309836 3856 309842 3868
rect 313936 3856 313964 3896
rect 325602 3884 325608 3896
rect 325660 3884 325666 3936
rect 327276 3896 329328 3924
rect 309836 3828 313964 3856
rect 314013 3859 314071 3865
rect 309836 3816 309842 3828
rect 314013 3825 314025 3859
rect 314059 3856 314071 3859
rect 326798 3856 326804 3868
rect 314059 3828 326804 3856
rect 314059 3825 314071 3828
rect 314013 3819 314071 3825
rect 326798 3816 326804 3828
rect 326856 3816 326862 3868
rect 258046 3760 258212 3788
rect 176654 3680 176660 3732
rect 176712 3720 176718 3732
rect 200758 3720 200764 3732
rect 176712 3692 200764 3720
rect 176712 3680 176718 3692
rect 200758 3680 200764 3692
rect 200816 3680 200822 3732
rect 229830 3680 229836 3732
rect 229888 3720 229894 3732
rect 258046 3720 258074 3760
rect 263042 3748 263048 3800
rect 263100 3788 263106 3800
rect 280338 3788 280344 3800
rect 263100 3760 280344 3788
rect 263100 3748 263106 3760
rect 280338 3748 280344 3760
rect 280396 3748 280402 3800
rect 304902 3748 304908 3800
rect 304960 3788 304966 3800
rect 318518 3788 318524 3800
rect 304960 3760 318524 3788
rect 304960 3748 304966 3760
rect 318518 3748 318524 3760
rect 318576 3748 318582 3800
rect 318702 3748 318708 3800
rect 318760 3788 318766 3800
rect 327276 3788 327304 3896
rect 329190 3856 329196 3868
rect 318760 3760 327304 3788
rect 327368 3828 329196 3856
rect 318760 3748 318766 3760
rect 262858 3720 262864 3732
rect 229888 3692 258074 3720
rect 258184 3692 262864 3720
rect 229888 3680 229894 3692
rect 179414 3652 179420 3664
rect 175660 3624 179420 3652
rect 179414 3612 179420 3624
rect 179472 3612 179478 3664
rect 180242 3612 180248 3664
rect 180300 3652 180306 3664
rect 204898 3652 204904 3664
rect 180300 3624 204904 3652
rect 180300 3612 180306 3624
rect 204898 3612 204904 3624
rect 204956 3612 204962 3664
rect 212166 3612 212172 3664
rect 212224 3652 212230 3664
rect 220078 3652 220084 3664
rect 212224 3624 220084 3652
rect 212224 3612 212230 3624
rect 220078 3612 220084 3624
rect 220136 3612 220142 3664
rect 226334 3612 226340 3664
rect 226392 3652 226398 3664
rect 258184 3652 258212 3692
rect 262858 3680 262864 3692
rect 262916 3680 262922 3732
rect 308950 3680 308956 3732
rect 309008 3720 309014 3732
rect 309008 3692 309180 3720
rect 309008 3680 309014 3692
rect 226392 3624 258212 3652
rect 226392 3612 226398 3624
rect 258258 3612 258264 3664
rect 258316 3652 258322 3664
rect 258718 3652 258724 3664
rect 258316 3624 258724 3652
rect 258316 3612 258322 3624
rect 258718 3612 258724 3624
rect 258776 3612 258782 3664
rect 265342 3612 265348 3664
rect 265400 3652 265406 3664
rect 280798 3652 280804 3664
rect 265400 3624 280804 3652
rect 265400 3612 265406 3624
rect 280798 3612 280804 3624
rect 280856 3612 280862 3664
rect 284294 3612 284300 3664
rect 284352 3652 284358 3664
rect 285490 3652 285496 3664
rect 284352 3624 285496 3652
rect 284352 3612 284358 3624
rect 285490 3612 285496 3624
rect 285548 3612 285554 3664
rect 305638 3612 305644 3664
rect 305696 3652 305702 3664
rect 309042 3652 309048 3664
rect 305696 3624 309048 3652
rect 305696 3612 305702 3624
rect 309042 3612 309048 3624
rect 309100 3612 309106 3664
rect 309152 3652 309180 3692
rect 313182 3680 313188 3732
rect 313240 3720 313246 3732
rect 313240 3692 316034 3720
rect 313240 3680 313246 3692
rect 314013 3655 314071 3661
rect 314013 3652 314025 3655
rect 309152 3624 314025 3652
rect 314013 3621 314025 3624
rect 314059 3621 314071 3655
rect 316006 3652 316034 3692
rect 316678 3680 316684 3732
rect 316736 3720 316742 3732
rect 317509 3723 317567 3729
rect 317509 3720 317521 3723
rect 316736 3692 317521 3720
rect 316736 3680 316742 3692
rect 317509 3689 317521 3692
rect 317555 3689 317567 3723
rect 317509 3683 317567 3689
rect 320821 3723 320879 3729
rect 320821 3689 320833 3723
rect 320867 3720 320879 3723
rect 327368 3720 327396 3828
rect 329190 3816 329196 3828
rect 329248 3816 329254 3868
rect 329300 3788 329328 3896
rect 335262 3884 335268 3936
rect 335320 3924 335326 3936
rect 387150 3924 387156 3936
rect 335320 3896 387156 3924
rect 335320 3884 335326 3896
rect 387150 3884 387156 3896
rect 387208 3884 387214 3936
rect 401502 3884 401508 3936
rect 401560 3924 401566 3936
rect 539594 3924 539600 3936
rect 401560 3896 539600 3924
rect 401560 3884 401566 3896
rect 539594 3884 539600 3896
rect 539652 3884 539658 3936
rect 336642 3816 336648 3868
rect 336700 3856 336706 3868
rect 390646 3856 390652 3868
rect 336700 3828 390652 3856
rect 336700 3816 336706 3828
rect 390646 3816 390652 3828
rect 390704 3816 390710 3868
rect 406378 3816 406384 3868
rect 406436 3856 406442 3868
rect 546678 3856 546684 3868
rect 406436 3828 546684 3856
rect 406436 3816 406442 3828
rect 546678 3816 546684 3828
rect 546736 3816 546742 3868
rect 348050 3788 348056 3800
rect 329300 3760 348056 3788
rect 348050 3748 348056 3760
rect 348108 3748 348114 3800
rect 352558 3748 352564 3800
rect 352616 3788 352622 3800
rect 408402 3788 408408 3800
rect 352616 3760 408408 3788
rect 352616 3748 352622 3760
rect 408402 3748 408408 3760
rect 408460 3748 408466 3800
rect 409138 3748 409144 3800
rect 409196 3788 409202 3800
rect 553762 3788 553768 3800
rect 409196 3760 553768 3788
rect 409196 3748 409202 3760
rect 553762 3748 553768 3760
rect 553820 3748 553826 3800
rect 320867 3692 327396 3720
rect 320867 3689 320879 3692
rect 320821 3683 320879 3689
rect 327718 3680 327724 3732
rect 327776 3720 327782 3732
rect 330386 3720 330392 3732
rect 327776 3692 330392 3720
rect 327776 3680 327782 3692
rect 330386 3680 330392 3692
rect 330444 3680 330450 3732
rect 330478 3680 330484 3732
rect 330536 3720 330542 3732
rect 333882 3720 333888 3732
rect 330536 3692 333888 3720
rect 330536 3680 330542 3692
rect 333882 3680 333888 3692
rect 333940 3680 333946 3732
rect 342162 3680 342168 3732
rect 342220 3720 342226 3732
rect 401318 3720 401324 3732
rect 342220 3692 401324 3720
rect 342220 3680 342226 3692
rect 401318 3680 401324 3692
rect 401376 3680 401382 3732
rect 411162 3680 411168 3732
rect 411220 3720 411226 3732
rect 560846 3720 560852 3732
rect 411220 3692 560852 3720
rect 411220 3680 411226 3692
rect 560846 3680 560852 3692
rect 560904 3680 560910 3732
rect 337470 3652 337476 3664
rect 316006 3624 337476 3652
rect 314013 3615 314071 3621
rect 337470 3612 337476 3624
rect 337528 3612 337534 3664
rect 339402 3612 339408 3664
rect 339460 3652 339466 3664
rect 397730 3652 397736 3664
rect 339460 3624 397736 3652
rect 339460 3612 339466 3624
rect 397730 3612 397736 3624
rect 397788 3612 397794 3664
rect 568022 3652 568028 3664
rect 419184 3624 568028 3652
rect 15930 3544 15936 3596
rect 15988 3584 15994 3596
rect 172514 3584 172520 3596
rect 15988 3556 172520 3584
rect 15988 3544 15994 3556
rect 172514 3544 172520 3556
rect 172572 3544 172578 3596
rect 188522 3544 188528 3596
rect 188580 3584 188586 3596
rect 244918 3584 244924 3596
rect 188580 3556 244924 3584
rect 188580 3544 188586 3556
rect 244918 3544 244924 3556
rect 244976 3544 244982 3596
rect 251174 3544 251180 3596
rect 251232 3584 251238 3596
rect 273898 3584 273904 3596
rect 251232 3556 273904 3584
rect 251232 3544 251238 3556
rect 273898 3544 273904 3556
rect 273956 3544 273962 3596
rect 276014 3544 276020 3596
rect 276072 3584 276078 3596
rect 277302 3584 277308 3596
rect 276072 3556 277308 3584
rect 276072 3544 276078 3556
rect 277302 3544 277308 3556
rect 277360 3544 277366 3596
rect 279510 3544 279516 3596
rect 279568 3584 279574 3596
rect 286318 3584 286324 3596
rect 279568 3556 286324 3584
rect 279568 3544 279574 3556
rect 286318 3544 286324 3556
rect 286376 3544 286382 3596
rect 303522 3544 303528 3596
rect 303580 3584 303586 3596
rect 303580 3556 306374 3584
rect 303580 3544 303586 3556
rect 5258 3476 5264 3528
rect 5316 3516 5322 3528
rect 11698 3516 11704 3528
rect 5316 3488 11704 3516
rect 5316 3476 5322 3488
rect 11698 3476 11704 3488
rect 11756 3476 11762 3528
rect 13538 3476 13544 3528
rect 13596 3516 13602 3528
rect 14550 3516 14556 3528
rect 13596 3488 14556 3516
rect 13596 3476 13602 3488
rect 14550 3476 14556 3488
rect 14608 3476 14614 3528
rect 14734 3476 14740 3528
rect 14792 3516 14798 3528
rect 171318 3516 171324 3528
rect 14792 3488 171324 3516
rect 14792 3476 14798 3488
rect 171318 3476 171324 3488
rect 171376 3476 171382 3528
rect 179046 3476 179052 3528
rect 179104 3516 179110 3528
rect 180058 3516 180064 3528
rect 179104 3488 180064 3516
rect 179104 3476 179110 3488
rect 180058 3476 180064 3488
rect 180116 3476 180122 3528
rect 185578 3516 185584 3528
rect 180766 3488 185584 3516
rect 6454 3408 6460 3460
rect 6512 3448 6518 3460
rect 164789 3451 164847 3457
rect 164789 3448 164801 3451
rect 6512 3420 164801 3448
rect 6512 3408 6518 3420
rect 164789 3417 164801 3420
rect 164835 3417 164847 3451
rect 164789 3411 164847 3417
rect 164878 3408 164884 3460
rect 164936 3448 164942 3460
rect 165522 3448 165528 3460
rect 164936 3420 165528 3448
rect 164936 3408 164942 3420
rect 165522 3408 165528 3420
rect 165580 3408 165586 3460
rect 166074 3408 166080 3460
rect 166132 3448 166138 3460
rect 166902 3448 166908 3460
rect 166132 3420 166908 3448
rect 166132 3408 166138 3420
rect 166902 3408 166908 3420
rect 166960 3408 166966 3460
rect 168374 3408 168380 3460
rect 168432 3448 168438 3460
rect 169570 3448 169576 3460
rect 168432 3420 169576 3448
rect 168432 3408 168438 3420
rect 169570 3408 169576 3420
rect 169628 3408 169634 3460
rect 18230 3340 18236 3392
rect 18288 3380 18294 3392
rect 19242 3380 19248 3392
rect 18288 3352 19248 3380
rect 18288 3340 18294 3352
rect 19242 3340 19248 3352
rect 19300 3340 19306 3392
rect 27706 3340 27712 3392
rect 27764 3380 27770 3392
rect 28902 3380 28908 3392
rect 27764 3352 28908 3380
rect 27764 3340 27770 3352
rect 28902 3340 28908 3352
rect 28960 3340 28966 3392
rect 31294 3340 31300 3392
rect 31352 3380 31358 3392
rect 32398 3380 32404 3392
rect 31352 3352 32404 3380
rect 31352 3340 31358 3352
rect 32398 3340 32404 3352
rect 32456 3340 32462 3392
rect 34790 3340 34796 3392
rect 34848 3380 34854 3392
rect 35802 3380 35808 3392
rect 34848 3352 35808 3380
rect 34848 3340 34854 3352
rect 35802 3340 35808 3352
rect 35860 3340 35866 3392
rect 38378 3340 38384 3392
rect 38436 3380 38442 3392
rect 39298 3380 39304 3392
rect 38436 3352 39304 3380
rect 38436 3340 38442 3352
rect 39298 3340 39304 3352
rect 39356 3340 39362 3392
rect 41874 3340 41880 3392
rect 41932 3380 41938 3392
rect 43438 3380 43444 3392
rect 41932 3352 43444 3380
rect 41932 3340 41938 3352
rect 43438 3340 43444 3352
rect 43496 3340 43502 3392
rect 58618 3380 58624 3392
rect 45526 3352 58624 3380
rect 43070 3272 43076 3324
rect 43128 3312 43134 3324
rect 45526 3312 45554 3352
rect 58618 3340 58624 3352
rect 58676 3340 58682 3392
rect 71498 3340 71504 3392
rect 71556 3380 71562 3392
rect 180766 3380 180794 3488
rect 185578 3476 185584 3488
rect 185636 3476 185642 3528
rect 186130 3476 186136 3528
rect 186188 3516 186194 3528
rect 188338 3516 188344 3528
rect 186188 3488 188344 3516
rect 186188 3476 186194 3488
rect 188338 3476 188344 3488
rect 188396 3476 188402 3528
rect 240413 3519 240471 3525
rect 240413 3516 240425 3519
rect 188448 3488 240425 3516
rect 183738 3408 183744 3460
rect 183796 3448 183802 3460
rect 188448 3448 188476 3488
rect 240413 3485 240425 3488
rect 240459 3485 240471 3519
rect 240413 3479 240471 3485
rect 240502 3476 240508 3528
rect 240560 3516 240566 3528
rect 241422 3516 241428 3528
rect 240560 3488 241428 3516
rect 240560 3476 240566 3488
rect 241422 3476 241428 3488
rect 241480 3476 241486 3528
rect 246390 3476 246396 3528
rect 246448 3516 246454 3528
rect 246942 3516 246948 3528
rect 246448 3488 246948 3516
rect 246448 3476 246454 3488
rect 246942 3476 246948 3488
rect 247000 3476 247006 3528
rect 247586 3476 247592 3528
rect 247644 3516 247650 3528
rect 271138 3516 271144 3528
rect 247644 3488 271144 3516
rect 247644 3476 247650 3488
rect 271138 3476 271144 3488
rect 271196 3476 271202 3528
rect 271230 3476 271236 3528
rect 271288 3516 271294 3528
rect 271782 3516 271788 3528
rect 271288 3488 271788 3516
rect 271288 3476 271294 3488
rect 271782 3476 271788 3488
rect 271840 3476 271846 3528
rect 274818 3476 274824 3528
rect 274876 3516 274882 3528
rect 276658 3516 276664 3528
rect 274876 3488 276664 3516
rect 274876 3476 274882 3488
rect 276658 3476 276664 3488
rect 276716 3476 276722 3528
rect 277118 3476 277124 3528
rect 277176 3516 277182 3528
rect 284938 3516 284944 3528
rect 277176 3488 284944 3516
rect 277176 3476 277182 3488
rect 284938 3476 284944 3488
rect 284996 3476 285002 3528
rect 288986 3476 288992 3528
rect 289044 3516 289050 3528
rect 289722 3516 289728 3528
rect 289044 3488 289728 3516
rect 289044 3476 289050 3488
rect 289722 3476 289728 3488
rect 289780 3476 289786 3528
rect 291378 3476 291384 3528
rect 291436 3516 291442 3528
rect 292482 3516 292488 3528
rect 291436 3488 292488 3516
rect 291436 3476 291442 3488
rect 292482 3476 292488 3488
rect 292540 3476 292546 3528
rect 294046 3476 294052 3528
rect 294104 3516 294110 3528
rect 294874 3516 294880 3528
rect 294104 3488 294880 3516
rect 294104 3476 294110 3488
rect 294874 3476 294880 3488
rect 294932 3476 294938 3528
rect 300118 3476 300124 3528
rect 300176 3516 300182 3528
rect 304350 3516 304356 3528
rect 300176 3488 304356 3516
rect 300176 3476 300182 3488
rect 304350 3476 304356 3488
rect 304408 3476 304414 3528
rect 306346 3516 306374 3556
rect 307662 3544 307668 3596
rect 307720 3584 307726 3596
rect 322106 3584 322112 3596
rect 307720 3556 322112 3584
rect 307720 3544 307726 3556
rect 322106 3544 322112 3556
rect 322164 3544 322170 3596
rect 322750 3544 322756 3596
rect 322808 3584 322814 3596
rect 357710 3584 357716 3596
rect 322808 3556 357716 3584
rect 322808 3544 322814 3556
rect 357710 3544 357716 3556
rect 357768 3544 357774 3596
rect 358262 3544 358268 3596
rect 358320 3584 358326 3596
rect 359918 3584 359924 3596
rect 358320 3556 359924 3584
rect 358320 3544 358326 3556
rect 359918 3544 359924 3556
rect 359976 3544 359982 3596
rect 360013 3587 360071 3593
rect 360013 3553 360025 3587
rect 360059 3584 360071 3587
rect 418982 3584 418988 3596
rect 360059 3556 418988 3584
rect 360059 3553 360071 3556
rect 360013 3547 360071 3553
rect 418982 3544 418988 3556
rect 419040 3544 419046 3596
rect 315022 3516 315028 3528
rect 306346 3488 315028 3516
rect 315022 3476 315028 3488
rect 315080 3476 315086 3528
rect 317230 3476 317236 3528
rect 317288 3516 317294 3528
rect 317509 3519 317567 3525
rect 317288 3488 317460 3516
rect 317288 3476 317294 3488
rect 244274 3448 244280 3460
rect 183796 3420 188476 3448
rect 190426 3420 244280 3448
rect 183796 3408 183802 3420
rect 71556 3352 180794 3380
rect 71556 3340 71562 3352
rect 181438 3340 181444 3392
rect 181496 3380 181502 3392
rect 190426 3380 190454 3420
rect 244274 3408 244280 3420
rect 244332 3408 244338 3460
rect 249978 3408 249984 3460
rect 250036 3448 250042 3460
rect 251082 3448 251088 3460
rect 250036 3420 251088 3448
rect 250036 3408 250042 3420
rect 251082 3408 251088 3420
rect 251140 3408 251146 3460
rect 253201 3451 253259 3457
rect 253201 3417 253213 3451
rect 253247 3448 253259 3451
rect 258166 3448 258172 3460
rect 253247 3420 258172 3448
rect 253247 3417 253259 3420
rect 253201 3411 253259 3417
rect 258166 3408 258172 3420
rect 258224 3408 258230 3460
rect 258258 3408 258264 3460
rect 258316 3448 258322 3460
rect 259362 3448 259368 3460
rect 258316 3420 259368 3448
rect 258316 3408 258322 3420
rect 259362 3408 259368 3420
rect 259420 3408 259426 3460
rect 259454 3408 259460 3460
rect 259512 3448 259518 3460
rect 260558 3448 260564 3460
rect 259512 3420 260564 3448
rect 259512 3408 259518 3420
rect 260558 3408 260564 3420
rect 260616 3408 260622 3460
rect 261754 3408 261760 3460
rect 261812 3448 261818 3460
rect 262950 3448 262956 3460
rect 261812 3420 262956 3448
rect 261812 3408 261818 3420
rect 262950 3408 262956 3420
rect 263008 3408 263014 3460
rect 264146 3408 264152 3460
rect 264204 3448 264210 3460
rect 264882 3448 264888 3460
rect 264204 3420 264888 3448
rect 264204 3408 264210 3420
rect 264882 3408 264888 3420
rect 264940 3408 264946 3460
rect 266538 3408 266544 3460
rect 266596 3448 266602 3460
rect 267642 3448 267648 3460
rect 266596 3420 267648 3448
rect 266596 3408 266602 3420
rect 267642 3408 267648 3420
rect 267700 3408 267706 3460
rect 273622 3408 273628 3460
rect 273680 3448 273686 3460
rect 282178 3448 282184 3460
rect 273680 3420 282184 3448
rect 273680 3408 273686 3420
rect 282178 3408 282184 3420
rect 282236 3408 282242 3460
rect 296530 3408 296536 3460
rect 296588 3448 296594 3460
rect 299658 3448 299664 3460
rect 296588 3420 299664 3448
rect 296588 3408 296594 3420
rect 299658 3408 299664 3420
rect 299716 3408 299722 3460
rect 304810 3408 304816 3460
rect 304868 3448 304874 3460
rect 317322 3448 317328 3460
rect 304868 3420 317328 3448
rect 304868 3408 304874 3420
rect 317322 3408 317328 3420
rect 317380 3408 317386 3460
rect 317432 3448 317460 3488
rect 317509 3485 317521 3519
rect 317555 3516 317567 3519
rect 340966 3516 340972 3528
rect 317555 3488 340972 3516
rect 317555 3485 317567 3488
rect 317509 3479 317567 3485
rect 340966 3476 340972 3488
rect 341024 3476 341030 3528
rect 343542 3476 343548 3528
rect 343600 3516 343606 3528
rect 404814 3516 404820 3528
rect 343600 3488 404820 3516
rect 343600 3476 343606 3488
rect 404814 3476 404820 3488
rect 404872 3476 404878 3528
rect 414658 3476 414664 3528
rect 414716 3516 414722 3528
rect 415486 3516 415492 3528
rect 414716 3488 415492 3516
rect 414716 3476 414722 3488
rect 415486 3476 415492 3488
rect 415544 3476 415550 3528
rect 344554 3448 344560 3460
rect 317432 3420 344560 3448
rect 344554 3408 344560 3420
rect 344612 3408 344618 3460
rect 346302 3408 346308 3460
rect 346360 3448 346366 3460
rect 411898 3448 411904 3460
rect 346360 3420 411904 3448
rect 346360 3408 346366 3420
rect 411898 3408 411904 3420
rect 411956 3408 411962 3460
rect 413922 3408 413928 3460
rect 413980 3448 413986 3460
rect 419184 3448 419212 3624
rect 568022 3612 568028 3624
rect 568080 3612 568086 3664
rect 419258 3544 419264 3596
rect 419316 3584 419322 3596
rect 575106 3584 575112 3596
rect 419316 3556 575112 3584
rect 419316 3544 419322 3556
rect 575106 3544 575112 3556
rect 575164 3544 575170 3596
rect 420822 3476 420828 3528
rect 420880 3516 420886 3528
rect 583386 3516 583392 3528
rect 420880 3488 583392 3516
rect 420880 3476 420886 3488
rect 583386 3476 583392 3488
rect 583444 3476 583450 3528
rect 413980 3420 419212 3448
rect 413980 3408 413986 3420
rect 419442 3408 419448 3460
rect 419500 3448 419506 3460
rect 580994 3448 581000 3460
rect 419500 3420 581000 3448
rect 419500 3408 419506 3420
rect 580994 3408 581000 3420
rect 581052 3408 581058 3460
rect 181496 3352 190454 3380
rect 181496 3340 181502 3352
rect 206186 3340 206192 3392
rect 206244 3380 206250 3392
rect 206922 3380 206928 3392
rect 206244 3352 206928 3380
rect 206244 3340 206250 3352
rect 206922 3340 206928 3352
rect 206980 3340 206986 3392
rect 208578 3340 208584 3392
rect 208636 3380 208642 3392
rect 209682 3380 209688 3392
rect 208636 3352 209688 3380
rect 208636 3340 208642 3352
rect 209682 3340 209688 3352
rect 209740 3340 209746 3392
rect 209774 3340 209780 3392
rect 209832 3380 209838 3392
rect 210970 3380 210976 3392
rect 209832 3352 210976 3380
rect 209832 3340 209838 3352
rect 210970 3340 210976 3352
rect 211028 3340 211034 3392
rect 213362 3340 213368 3392
rect 213420 3380 213426 3392
rect 213822 3380 213828 3392
rect 213420 3352 213828 3380
rect 213420 3340 213426 3352
rect 213822 3340 213828 3352
rect 213880 3340 213886 3392
rect 215662 3340 215668 3392
rect 215720 3380 215726 3392
rect 216582 3380 216588 3392
rect 215720 3352 216588 3380
rect 215720 3340 215726 3352
rect 216582 3340 216588 3352
rect 216640 3340 216646 3392
rect 216858 3340 216864 3392
rect 216916 3380 216922 3392
rect 217962 3380 217968 3392
rect 216916 3352 217968 3380
rect 216916 3340 216922 3352
rect 217962 3340 217968 3352
rect 218020 3340 218026 3392
rect 222746 3340 222752 3392
rect 222804 3380 222810 3392
rect 223482 3380 223488 3392
rect 222804 3352 223488 3380
rect 222804 3340 222810 3352
rect 223482 3340 223488 3352
rect 223540 3340 223546 3392
rect 231026 3340 231032 3392
rect 231084 3380 231090 3392
rect 231762 3380 231768 3392
rect 231084 3352 231768 3380
rect 231084 3340 231090 3352
rect 231762 3340 231768 3352
rect 231820 3340 231826 3392
rect 233418 3340 233424 3392
rect 233476 3380 233482 3392
rect 234522 3380 234528 3392
rect 233476 3352 234528 3380
rect 233476 3340 233482 3352
rect 234522 3340 234528 3352
rect 234580 3340 234586 3392
rect 235810 3340 235816 3392
rect 235868 3380 235874 3392
rect 240413 3383 240471 3389
rect 235868 3352 240364 3380
rect 235868 3340 235874 3352
rect 43128 3284 45554 3312
rect 43128 3272 43134 3284
rect 60826 3272 60832 3324
rect 60884 3312 60890 3324
rect 71038 3312 71044 3324
rect 60884 3284 71044 3312
rect 60884 3272 60890 3284
rect 71038 3272 71044 3284
rect 71096 3272 71102 3324
rect 78582 3272 78588 3324
rect 78640 3312 78646 3324
rect 186958 3312 186964 3324
rect 78640 3284 186964 3312
rect 78640 3272 78646 3284
rect 186958 3272 186964 3284
rect 187016 3272 187022 3324
rect 234614 3272 234620 3324
rect 234672 3312 234678 3324
rect 235902 3312 235908 3324
rect 234672 3284 235908 3312
rect 234672 3272 234678 3284
rect 235902 3272 235908 3284
rect 235960 3272 235966 3324
rect 238110 3272 238116 3324
rect 238168 3312 238174 3324
rect 238662 3312 238668 3324
rect 238168 3284 238668 3312
rect 238168 3272 238174 3284
rect 238662 3272 238668 3284
rect 238720 3272 238726 3324
rect 240336 3312 240364 3352
rect 240413 3349 240425 3383
rect 240459 3380 240471 3383
rect 245838 3380 245844 3392
rect 240459 3352 245844 3380
rect 240459 3349 240471 3352
rect 240413 3343 240471 3349
rect 245838 3340 245844 3352
rect 245896 3340 245902 3392
rect 254670 3340 254676 3392
rect 254728 3380 254734 3392
rect 254728 3352 272012 3380
rect 254728 3340 254734 3352
rect 245010 3312 245016 3324
rect 240336 3284 245016 3312
rect 245010 3272 245016 3284
rect 245068 3272 245074 3324
rect 245194 3272 245200 3324
rect 245252 3312 245258 3324
rect 251818 3312 251824 3324
rect 245252 3284 251824 3312
rect 245252 3272 245258 3284
rect 251818 3272 251824 3284
rect 251876 3272 251882 3324
rect 255866 3272 255872 3324
rect 255924 3312 255930 3324
rect 271984 3312 272012 3352
rect 272426 3340 272432 3392
rect 272484 3380 272490 3392
rect 282270 3380 282276 3392
rect 272484 3352 282276 3380
rect 272484 3340 272490 3352
rect 282270 3340 282276 3352
rect 282328 3340 282334 3392
rect 304258 3340 304264 3392
rect 304316 3380 304322 3392
rect 311434 3380 311440 3392
rect 304316 3352 311440 3380
rect 304316 3340 304322 3352
rect 311434 3340 311440 3352
rect 311492 3340 311498 3392
rect 324222 3340 324228 3392
rect 324280 3380 324286 3392
rect 361114 3380 361120 3392
rect 324280 3352 361120 3380
rect 324280 3340 324286 3352
rect 361114 3340 361120 3352
rect 361172 3340 361178 3392
rect 363598 3340 363604 3392
rect 363656 3380 363662 3392
rect 447410 3380 447416 3392
rect 363656 3352 447416 3380
rect 363656 3340 363662 3352
rect 447410 3340 447416 3352
rect 447468 3340 447474 3392
rect 448514 3340 448520 3392
rect 448572 3380 448578 3392
rect 449802 3380 449808 3392
rect 448572 3352 449808 3380
rect 448572 3340 448578 3352
rect 449802 3340 449808 3352
rect 449860 3340 449866 3392
rect 456794 3340 456800 3392
rect 456852 3380 456858 3392
rect 458082 3380 458088 3392
rect 456852 3352 458088 3380
rect 456852 3340 456858 3352
rect 458082 3340 458088 3352
rect 458140 3340 458146 3392
rect 482186 3340 482192 3392
rect 482244 3380 482250 3392
rect 571518 3380 571524 3392
rect 482244 3352 571524 3380
rect 482244 3340 482250 3352
rect 571518 3340 571524 3352
rect 571576 3340 571582 3392
rect 276198 3312 276204 3324
rect 255924 3284 267734 3312
rect 271984 3284 276204 3312
rect 255924 3272 255930 3284
rect 9950 3204 9956 3256
rect 10008 3244 10014 3256
rect 14458 3244 14464 3256
rect 10008 3216 14464 3244
rect 10008 3204 10014 3216
rect 14458 3204 14464 3216
rect 14516 3204 14522 3256
rect 28902 3204 28908 3256
rect 28960 3244 28966 3256
rect 35158 3244 35164 3256
rect 28960 3216 35164 3244
rect 28960 3204 28966 3216
rect 35158 3204 35164 3216
rect 35216 3204 35222 3256
rect 89162 3204 89168 3256
rect 89220 3244 89226 3256
rect 189626 3244 189632 3256
rect 89220 3216 189632 3244
rect 89220 3204 89226 3216
rect 189626 3204 189632 3216
rect 189684 3204 189690 3256
rect 239306 3204 239312 3256
rect 239364 3244 239370 3256
rect 260098 3244 260104 3256
rect 239364 3216 260104 3244
rect 239364 3204 239370 3216
rect 260098 3204 260104 3216
rect 260156 3204 260162 3256
rect 267706 3244 267734 3284
rect 276198 3272 276204 3284
rect 276256 3272 276262 3324
rect 280706 3272 280712 3324
rect 280764 3312 280770 3324
rect 287330 3312 287336 3324
rect 280764 3284 287336 3312
rect 280764 3272 280770 3284
rect 287330 3272 287336 3284
rect 287388 3272 287394 3324
rect 310422 3272 310428 3324
rect 310480 3312 310486 3324
rect 320821 3315 320879 3321
rect 320821 3312 320833 3315
rect 310480 3284 320833 3312
rect 310480 3272 310486 3284
rect 320821 3281 320833 3284
rect 320867 3281 320879 3315
rect 320821 3275 320879 3281
rect 325418 3272 325424 3324
rect 325476 3312 325482 3324
rect 365806 3312 365812 3324
rect 325476 3284 365812 3312
rect 325476 3272 325482 3284
rect 365806 3272 365812 3284
rect 365864 3272 365870 3324
rect 368937 3315 368995 3321
rect 368937 3281 368949 3315
rect 368983 3312 368995 3315
rect 376478 3312 376484 3324
rect 368983 3284 376484 3312
rect 368983 3281 368995 3284
rect 368937 3275 368995 3281
rect 376478 3272 376484 3284
rect 376536 3272 376542 3324
rect 378778 3272 378784 3324
rect 378836 3312 378842 3324
rect 461578 3312 461584 3324
rect 378836 3284 461584 3312
rect 378836 3272 378842 3284
rect 461578 3272 461584 3284
rect 461636 3272 461642 3324
rect 479518 3272 479524 3324
rect 479576 3312 479582 3324
rect 564434 3312 564440 3324
rect 479576 3284 564440 3312
rect 479576 3272 479582 3284
rect 564434 3272 564440 3284
rect 564492 3272 564498 3324
rect 277578 3244 277584 3256
rect 267706 3216 277584 3244
rect 277578 3204 277584 3216
rect 277636 3204 277642 3256
rect 325510 3204 325516 3256
rect 325568 3244 325574 3256
rect 364610 3244 364616 3256
rect 325568 3216 364616 3244
rect 325568 3204 325574 3216
rect 364610 3204 364616 3216
rect 364668 3204 364674 3256
rect 376018 3204 376024 3256
rect 376076 3244 376082 3256
rect 454494 3244 454500 3256
rect 376076 3216 454500 3244
rect 376076 3204 376082 3216
rect 454494 3204 454500 3216
rect 454552 3204 454558 3256
rect 478230 3204 478236 3256
rect 478288 3244 478294 3256
rect 557350 3244 557356 3256
rect 478288 3216 557356 3244
rect 478288 3204 478294 3216
rect 557350 3204 557356 3216
rect 557408 3204 557414 3256
rect 96246 3136 96252 3188
rect 96304 3176 96310 3188
rect 191098 3176 191104 3188
rect 96304 3148 191104 3176
rect 96304 3136 96310 3148
rect 191098 3136 191104 3148
rect 191156 3136 191162 3188
rect 257062 3136 257068 3188
rect 257120 3176 257126 3188
rect 268378 3176 268384 3188
rect 257120 3148 268384 3176
rect 257120 3136 257126 3148
rect 268378 3136 268384 3148
rect 268436 3136 268442 3188
rect 287790 3136 287796 3188
rect 287848 3176 287854 3188
rect 291286 3176 291292 3188
rect 287848 3148 291292 3176
rect 287848 3136 287854 3148
rect 291286 3136 291292 3148
rect 291344 3136 291350 3188
rect 298738 3136 298744 3188
rect 298796 3176 298802 3188
rect 301958 3176 301964 3188
rect 298796 3148 301964 3176
rect 298796 3136 298802 3148
rect 301958 3136 301964 3148
rect 302016 3136 302022 3188
rect 307018 3136 307024 3188
rect 307076 3176 307082 3188
rect 310238 3176 310244 3188
rect 307076 3148 310244 3176
rect 307076 3136 307082 3148
rect 310238 3136 310244 3148
rect 310296 3136 310302 3188
rect 322842 3136 322848 3188
rect 322900 3176 322906 3188
rect 357526 3176 357532 3188
rect 322900 3148 357532 3176
rect 322900 3136 322906 3148
rect 357526 3136 357532 3148
rect 357584 3136 357590 3188
rect 358170 3136 358176 3188
rect 358228 3176 358234 3188
rect 360013 3179 360071 3185
rect 360013 3176 360025 3179
rect 358228 3148 360025 3176
rect 358228 3136 358234 3148
rect 360013 3145 360025 3148
rect 360059 3145 360071 3179
rect 360013 3139 360071 3145
rect 360930 3136 360936 3188
rect 360988 3176 360994 3188
rect 360988 3148 364334 3176
rect 360988 3136 360994 3148
rect 74994 3068 75000 3120
rect 75052 3108 75058 3120
rect 98546 3108 98552 3120
rect 75052 3080 98552 3108
rect 75052 3068 75058 3080
rect 98546 3068 98552 3080
rect 98604 3068 98610 3120
rect 103330 3068 103336 3120
rect 103388 3108 103394 3120
rect 192478 3108 192484 3120
rect 103388 3080 192484 3108
rect 103388 3068 103394 3080
rect 192478 3068 192484 3080
rect 192536 3068 192542 3120
rect 248782 3068 248788 3120
rect 248840 3108 248846 3120
rect 273438 3108 273444 3120
rect 248840 3080 273444 3108
rect 248840 3068 248846 3080
rect 273438 3068 273444 3080
rect 273496 3068 273502 3120
rect 283098 3068 283104 3120
rect 283156 3108 283162 3120
rect 287698 3108 287704 3120
rect 283156 3080 287704 3108
rect 283156 3068 283162 3080
rect 287698 3068 287704 3080
rect 287756 3068 287762 3120
rect 321370 3068 321376 3120
rect 321428 3108 321434 3120
rect 355226 3108 355232 3120
rect 321428 3080 355232 3108
rect 321428 3068 321434 3080
rect 355226 3068 355232 3080
rect 355284 3068 355290 3120
rect 356698 3068 356704 3120
rect 356756 3108 356762 3120
rect 362310 3108 362316 3120
rect 356756 3080 362316 3108
rect 356756 3068 356762 3080
rect 362310 3068 362316 3080
rect 362368 3068 362374 3120
rect 364306 3108 364334 3148
rect 364978 3136 364984 3188
rect 365036 3176 365042 3188
rect 440326 3176 440332 3188
rect 365036 3148 440332 3176
rect 365036 3136 365042 3148
rect 440326 3136 440332 3148
rect 440384 3136 440390 3188
rect 473998 3136 474004 3188
rect 474056 3176 474062 3188
rect 550266 3176 550272 3188
rect 474056 3148 550272 3176
rect 474056 3136 474062 3148
rect 550266 3136 550272 3148
rect 550324 3136 550330 3188
rect 383562 3108 383568 3120
rect 364306 3080 383568 3108
rect 383562 3068 383568 3080
rect 383620 3068 383626 3120
rect 393958 3068 393964 3120
rect 394016 3108 394022 3120
rect 465166 3108 465172 3120
rect 394016 3080 465172 3108
rect 394016 3068 394022 3080
rect 465166 3068 465172 3080
rect 465224 3068 465230 3120
rect 472618 3068 472624 3120
rect 472676 3108 472682 3120
rect 543182 3108 543188 3120
rect 472676 3080 543188 3108
rect 472676 3068 472682 3080
rect 543182 3068 543188 3080
rect 543240 3068 543246 3120
rect 82078 3000 82084 3052
rect 82136 3040 82142 3052
rect 105538 3040 105544 3052
rect 82136 3012 105544 3040
rect 82136 3000 82142 3012
rect 105538 3000 105544 3012
rect 105596 3000 105602 3052
rect 110506 3000 110512 3052
rect 110564 3040 110570 3052
rect 193858 3040 193864 3052
rect 110564 3012 193864 3040
rect 110564 3000 110570 3012
rect 193858 3000 193864 3012
rect 193916 3000 193922 3052
rect 252370 3000 252376 3052
rect 252428 3040 252434 3052
rect 255958 3040 255964 3052
rect 252428 3012 255964 3040
rect 252428 3000 252434 3012
rect 255958 3000 255964 3012
rect 256016 3000 256022 3052
rect 298830 3000 298836 3052
rect 298888 3040 298894 3052
rect 300762 3040 300768 3052
rect 298888 3012 300768 3040
rect 298888 3000 298894 3012
rect 300762 3000 300768 3012
rect 300820 3000 300826 3052
rect 321462 3000 321468 3052
rect 321520 3040 321526 3052
rect 354030 3040 354036 3052
rect 321520 3012 354036 3040
rect 321520 3000 321526 3012
rect 354030 3000 354036 3012
rect 354088 3000 354094 3052
rect 360838 3000 360844 3052
rect 360896 3040 360902 3052
rect 433242 3040 433248 3052
rect 360896 3012 433248 3040
rect 360896 3000 360902 3012
rect 433242 3000 433248 3012
rect 433300 3000 433306 3052
rect 471238 3000 471244 3052
rect 471296 3040 471302 3052
rect 536098 3040 536104 3052
rect 471296 3012 536104 3040
rect 471296 3000 471302 3012
rect 536098 3000 536104 3012
rect 536156 3000 536162 3052
rect 85666 2932 85672 2984
rect 85724 2972 85730 2984
rect 111058 2972 111064 2984
rect 85724 2944 111064 2972
rect 85724 2932 85730 2944
rect 111058 2932 111064 2944
rect 111116 2932 111122 2984
rect 117590 2932 117596 2984
rect 117648 2972 117654 2984
rect 195238 2972 195244 2984
rect 117648 2944 195244 2972
rect 117648 2932 117654 2944
rect 195238 2932 195244 2944
rect 195296 2932 195302 2984
rect 195606 2932 195612 2984
rect 195664 2972 195670 2984
rect 198090 2972 198096 2984
rect 195664 2944 198096 2972
rect 195664 2932 195670 2944
rect 198090 2932 198096 2944
rect 198148 2932 198154 2984
rect 290182 2932 290188 2984
rect 290240 2972 290246 2984
rect 291470 2972 291476 2984
rect 290240 2944 291476 2972
rect 290240 2932 290246 2944
rect 291470 2932 291476 2944
rect 291528 2932 291534 2984
rect 322198 2932 322204 2984
rect 322256 2972 322262 2984
rect 351638 2972 351644 2984
rect 322256 2944 351644 2972
rect 322256 2932 322262 2944
rect 351638 2932 351644 2944
rect 351696 2932 351702 2984
rect 359458 2932 359464 2984
rect 359516 2972 359522 2984
rect 426158 2972 426164 2984
rect 359516 2944 426164 2972
rect 359516 2932 359522 2944
rect 426158 2932 426164 2944
rect 426216 2932 426222 2984
rect 467190 2932 467196 2984
rect 467248 2972 467254 2984
rect 467248 2944 509234 2972
rect 467248 2932 467254 2944
rect 121086 2864 121092 2916
rect 121144 2904 121150 2916
rect 196618 2904 196624 2916
rect 121144 2876 196624 2904
rect 121144 2864 121150 2876
rect 196618 2864 196624 2876
rect 196676 2864 196682 2916
rect 267734 2864 267740 2916
rect 267792 2904 267798 2916
rect 269022 2904 269028 2916
rect 267792 2876 269028 2904
rect 267792 2864 267798 2876
rect 269022 2864 269028 2876
rect 269080 2864 269086 2916
rect 335998 2864 336004 2916
rect 336056 2904 336062 2916
rect 350442 2904 350448 2916
rect 336056 2876 350448 2904
rect 336056 2864 336062 2876
rect 350442 2864 350448 2876
rect 350500 2864 350506 2916
rect 353938 2864 353944 2916
rect 353996 2904 354002 2916
rect 368198 2904 368204 2916
rect 353996 2876 368204 2904
rect 353996 2864 354002 2876
rect 368198 2864 368204 2876
rect 368256 2864 368262 2916
rect 509206 2904 509234 2944
rect 522298 2932 522304 2984
rect 522356 2972 522362 2984
rect 524230 2972 524236 2984
rect 522356 2944 524236 2972
rect 522356 2932 522362 2944
rect 524230 2932 524236 2944
rect 524288 2932 524294 2984
rect 529014 2904 529020 2916
rect 509206 2876 529020 2904
rect 529014 2864 529020 2876
rect 529072 2864 529078 2916
rect 25314 2796 25320 2848
rect 25372 2836 25378 2848
rect 176838 2836 176844 2848
rect 25372 2808 176844 2836
rect 25372 2796 25378 2808
rect 176838 2796 176844 2808
rect 176896 2796 176902 2848
rect 182542 2796 182548 2848
rect 182600 2836 182606 2848
rect 196710 2836 196716 2848
rect 182600 2808 196716 2836
rect 182600 2796 182606 2808
rect 196710 2796 196716 2808
rect 196768 2796 196774 2848
rect 357710 2796 357716 2848
rect 357768 2836 357774 2848
rect 358722 2836 358728 2848
rect 357768 2808 358728 2836
rect 357768 2796 357774 2808
rect 358722 2796 358728 2808
rect 358780 2796 358786 2848
rect 359550 2796 359556 2848
rect 359608 2836 359614 2848
rect 369394 2836 369400 2848
rect 359608 2808 369400 2836
rect 359608 2796 359614 2808
rect 369394 2796 369400 2808
rect 369452 2796 369458 2848
<< via1 >>
rect 137836 700952 137888 701004
rect 309140 700952 309192 701004
rect 277308 700884 277360 700936
rect 462320 700884 462372 700936
rect 278688 700816 278740 700868
rect 478512 700816 478564 700868
rect 105452 700748 105504 700800
rect 313280 700748 313332 700800
rect 89168 700680 89220 700732
rect 317420 700680 317472 700732
rect 72976 700612 73028 700664
rect 316040 700612 316092 700664
rect 270408 700544 270460 700596
rect 527180 700544 527232 700596
rect 271788 700476 271840 700528
rect 543464 700476 543516 700528
rect 40500 700408 40552 700460
rect 320180 700408 320232 700460
rect 24308 700340 24360 700392
rect 324320 700340 324372 700392
rect 8116 700272 8168 700324
rect 322940 700272 322992 700324
rect 154120 700204 154172 700256
rect 311900 700204 311952 700256
rect 285588 700136 285640 700188
rect 413652 700136 413704 700188
rect 202788 700068 202840 700120
rect 302240 700068 302292 700120
rect 302884 700068 302936 700120
rect 429844 700068 429896 700120
rect 284208 700000 284260 700052
rect 397460 700000 397512 700052
rect 292488 699932 292540 699984
rect 348792 699932 348844 699984
rect 289728 699864 289780 699916
rect 332508 699864 332560 699916
rect 267648 699796 267700 699848
rect 295340 699796 295392 699848
rect 283840 699728 283892 699780
rect 298100 699728 298152 699780
rect 170312 699660 170364 699712
rect 171048 699660 171100 699712
rect 235172 699660 235224 699712
rect 235908 699660 235960 699712
rect 263508 696940 263560 696992
rect 580172 696940 580224 696992
rect 266268 683204 266320 683256
rect 580172 683204 580224 683256
rect 3424 683136 3476 683188
rect 327080 683136 327132 683188
rect 260748 670760 260800 670812
rect 580172 670760 580224 670812
rect 3516 670692 3568 670744
rect 331220 670692 331272 670744
rect 3424 656888 3476 656940
rect 329840 656888 329892 656940
rect 256608 643084 256660 643136
rect 580172 643084 580224 643136
rect 3424 632068 3476 632120
rect 333980 632068 334032 632120
rect 259368 630640 259420 630692
rect 580172 630640 580224 630692
rect 3148 618264 3200 618316
rect 338120 618264 338172 618316
rect 255228 616836 255280 616888
rect 580172 616836 580224 616888
rect 3240 605820 3292 605872
rect 335360 605820 335412 605872
rect 249708 590656 249760 590708
rect 579804 590656 579856 590708
rect 3332 579640 3384 579692
rect 340880 579640 340932 579692
rect 252468 576852 252520 576904
rect 580172 576852 580224 576904
rect 3424 565836 3476 565888
rect 345020 565836 345072 565888
rect 248328 563048 248380 563100
rect 579804 563048 579856 563100
rect 3424 553392 3476 553444
rect 342260 553392 342312 553444
rect 242808 536800 242860 536852
rect 580172 536800 580224 536852
rect 3424 527144 3476 527196
rect 347780 527144 347832 527196
rect 245568 524424 245620 524476
rect 580172 524424 580224 524476
rect 3424 514768 3476 514820
rect 351920 514768 351972 514820
rect 294144 511708 294196 511760
rect 299480 511708 299532 511760
rect 280712 511640 280764 511692
rect 302884 511640 302936 511692
rect 235908 511572 235960 511624
rect 300860 511572 300912 511624
rect 287428 511504 287480 511556
rect 364340 511504 364392 511556
rect 219348 511436 219400 511488
rect 305276 511436 305328 511488
rect 171048 511368 171100 511420
rect 307576 511368 307628 511420
rect 274088 511300 274140 511352
rect 494060 511300 494112 511352
rect 267372 511232 267424 511284
rect 558920 511232 558972 511284
rect 240508 510620 240560 510672
rect 580172 510620 580224 510672
rect 198096 510552 198148 510604
rect 237380 510552 237432 510604
rect 238300 510552 238352 510604
rect 431316 510552 431368 510604
rect 231584 510484 231636 510536
rect 431224 510484 431276 510536
rect 229376 510416 229428 510468
rect 430120 510416 430172 510468
rect 175832 510348 175884 510400
rect 424324 510348 424376 510400
rect 215944 510280 215996 510332
rect 478144 510280 478196 510332
rect 224960 510212 225012 510264
rect 496084 510212 496136 510264
rect 100116 510144 100168 510196
rect 399116 510144 399168 510196
rect 101496 510076 101548 510128
rect 405832 510076 405884 510128
rect 100024 510008 100076 510060
rect 412456 510008 412508 510060
rect 101404 509940 101456 509992
rect 419172 509940 419224 509992
rect 82084 509872 82136 509924
rect 410248 509872 410300 509924
rect 64144 509804 64196 509856
rect 403532 509804 403584 509856
rect 222660 509736 222712 509788
rect 562324 509736 562376 509788
rect 4988 509668 5040 509720
rect 365628 509668 365680 509720
rect 14648 509600 14700 509652
rect 376760 509600 376812 509652
rect 4896 509532 4948 509584
rect 372344 509532 372396 509584
rect 11704 509464 11756 509516
rect 378968 509464 379020 509516
rect 14556 509396 14608 509448
rect 385684 509396 385736 509448
rect 14464 509328 14516 509380
rect 392400 509328 392452 509380
rect 4804 509260 4856 509312
rect 390192 509260 390244 509312
rect 237380 509235 237432 509244
rect 237380 509201 237389 509235
rect 237389 509201 237423 509235
rect 237423 509201 237432 509235
rect 237380 509192 237432 509201
rect 233884 509124 233936 509176
rect 421932 509124 421984 509176
rect 213736 509056 213788 509108
rect 425888 509056 425940 509108
rect 207020 508988 207072 509040
rect 424508 508988 424560 509040
rect 200396 508920 200448 508972
rect 422944 508920 422996 508972
rect 193680 508852 193732 508904
rect 424416 508852 424468 508904
rect 186964 508784 187016 508836
rect 421840 508784 421892 508836
rect 180248 508716 180300 508768
rect 421748 508716 421800 508768
rect 173532 508648 173584 508700
rect 421656 508648 421708 508700
rect 169116 508580 169168 508632
rect 508504 508580 508556 508632
rect 7932 508512 7984 508564
rect 354404 508512 354456 508564
rect 7840 508444 7892 508496
rect 361120 508512 361172 508564
rect 356704 508487 356756 508496
rect 356704 508453 356713 508487
rect 356713 508453 356747 508487
rect 356747 508453 356756 508487
rect 356704 508444 356756 508453
rect 358912 508487 358964 508496
rect 358912 508453 358921 508487
rect 358921 508453 358955 508487
rect 358955 508453 358964 508487
rect 358912 508444 358964 508453
rect 363328 508487 363380 508496
rect 363328 508453 363337 508487
rect 363337 508453 363371 508487
rect 363371 508453 363380 508487
rect 363328 508444 363380 508453
rect 220452 508376 220504 508428
rect 573364 508376 573416 508428
rect 7748 508308 7800 508360
rect 367836 508308 367888 508360
rect 370044 508351 370096 508360
rect 370044 508317 370053 508351
rect 370053 508317 370087 508351
rect 370087 508317 370096 508351
rect 370044 508308 370096 508317
rect 9036 508240 9088 508292
rect 374552 508240 374604 508292
rect 10508 508172 10560 508224
rect 381268 508172 381320 508224
rect 383476 508215 383528 508224
rect 383476 508181 383485 508215
rect 383485 508181 383519 508215
rect 383519 508181 383528 508215
rect 383476 508172 383528 508181
rect 8944 508104 8996 508156
rect 387892 508104 387944 508156
rect 10416 508036 10468 508088
rect 394608 508036 394660 508088
rect 7656 507968 7708 508020
rect 401324 508036 401376 508088
rect 396540 508011 396592 508020
rect 396540 507977 396549 508011
rect 396549 507977 396583 508011
rect 396583 507977 396592 508011
rect 396540 507968 396592 507977
rect 7564 507900 7616 507952
rect 407764 507900 407816 507952
rect 10324 507832 10376 507884
rect 414388 507832 414440 507884
rect 236368 507764 236420 507816
rect 426072 507764 426124 507816
rect 211896 507696 211948 507748
rect 218520 507671 218572 507680
rect 218520 507637 218529 507671
rect 218529 507637 218563 507671
rect 218563 507637 218572 507671
rect 218520 507628 218572 507637
rect 227536 507696 227588 507748
rect 425980 507696 426032 507748
rect 429936 507628 429988 507680
rect 205088 507603 205140 507612
rect 205088 507569 205097 507603
rect 205097 507569 205131 507603
rect 205131 507569 205140 507603
rect 205088 507560 205140 507569
rect 209504 507560 209556 507612
rect 430028 507560 430080 507612
rect 202788 507492 202840 507544
rect 428740 507492 428792 507544
rect 195796 507424 195848 507476
rect 428648 507424 428700 507476
rect 191656 507356 191708 507408
rect 429844 507356 429896 507408
rect 182824 507288 182876 507340
rect 184940 507220 184992 507272
rect 189448 507288 189500 507340
rect 428556 507288 428608 507340
rect 349712 507220 349764 507272
rect 425796 507220 425848 507272
rect 5540 507016 5592 507068
rect 428464 507152 428516 507204
rect 580264 507084 580316 507136
rect 11980 506948 12032 507000
rect 11888 506880 11940 506932
rect 5080 506812 5132 506864
rect 11796 506744 11848 506796
rect 580448 506676 580500 506728
rect 580356 506608 580408 506660
rect 3608 506540 3660 506592
rect 3516 506472 3568 506524
rect 3148 502256 3200 502308
rect 5540 502256 5592 502308
rect 426072 485732 426124 485784
rect 580172 485732 580224 485784
rect 3332 475668 3384 475720
rect 7932 475668 7984 475720
rect 431316 471928 431368 471980
rect 580172 471928 580224 471980
rect 2780 463428 2832 463480
rect 5080 463428 5132 463480
rect 421932 458124 421984 458176
rect 580172 458124 580224 458176
rect 3332 449828 3384 449880
rect 11980 449828 12032 449880
rect 430120 431876 430172 431928
rect 580172 431876 580224 431928
rect 3332 423580 3384 423632
rect 7840 423580 7892 423632
rect 431224 419432 431276 419484
rect 579712 419432 579764 419484
rect 2780 411000 2832 411052
rect 4988 411000 5040 411052
rect 425980 405628 426032 405680
rect 579804 405628 579856 405680
rect 3332 398760 3384 398812
rect 11888 398760 11940 398812
rect 562324 379448 562376 379500
rect 579804 379448 579856 379500
rect 3056 372376 3108 372428
rect 7748 372376 7800 372428
rect 496084 365644 496136 365696
rect 580172 365644 580224 365696
rect 2780 358436 2832 358488
rect 4896 358436 4948 358488
rect 573364 353200 573416 353252
rect 579620 353200 579672 353252
rect 3332 346332 3384 346384
rect 11796 346332 11848 346384
rect 478144 325592 478196 325644
rect 580172 325592 580224 325644
rect 3332 319540 3384 319592
rect 9036 319540 9088 319592
rect 3332 306280 3384 306332
rect 11704 306280 11756 306332
rect 425888 299412 425940 299464
rect 580172 299412 580224 299464
rect 2872 293904 2924 293956
rect 14648 293904 14700 293956
rect 430028 273164 430080 273216
rect 580172 273164 580224 273216
rect 3240 267656 3292 267708
rect 10508 267656 10560 267708
rect 429936 259360 429988 259412
rect 579620 259360 579672 259412
rect 3332 255212 3384 255264
rect 14556 255212 14608 255264
rect 424508 245556 424560 245608
rect 580172 245556 580224 245608
rect 428740 233180 428792 233232
rect 580172 233180 580224 233232
rect 3332 214956 3384 215008
rect 8944 214956 8996 215008
rect 422944 206932 422996 206984
rect 580172 206932 580224 206984
rect 3056 202784 3108 202836
rect 14464 202784 14516 202836
rect 168472 200404 168524 200456
rect 168748 200404 168800 200456
rect 240232 200404 240284 200456
rect 240508 200404 240560 200456
rect 252560 200404 252612 200456
rect 252836 200404 252888 200456
rect 61384 198636 61436 198688
rect 174452 198636 174504 198688
rect 177304 198636 177356 198688
rect 218152 198636 218204 198688
rect 238668 198636 238720 198688
rect 269396 198636 269448 198688
rect 277308 198636 277360 198688
rect 285956 198636 286008 198688
rect 312912 198636 312964 198688
rect 335544 198636 335596 198688
rect 337936 198636 337988 198688
rect 393504 198636 393556 198688
rect 395528 198636 395580 198688
rect 400128 198636 400180 198688
rect 471244 198636 471296 198688
rect 76564 198568 76616 198620
rect 195060 198568 195112 198620
rect 196900 198568 196952 198620
rect 213092 198568 213144 198620
rect 213276 198568 213328 198620
rect 229652 198568 229704 198620
rect 235908 198568 235960 198620
rect 267924 198568 267976 198620
rect 271788 198568 271840 198620
rect 283932 198568 283984 198620
rect 319168 198568 319220 198620
rect 336004 198568 336056 198620
rect 347504 198568 347556 198620
rect 414572 198568 414624 198620
rect 419356 198568 419408 198620
rect 490564 198568 490616 198620
rect 71044 198500 71096 198552
rect 191932 198500 191984 198552
rect 198004 198500 198056 198552
rect 214748 198500 214800 198552
rect 217324 198500 217376 198552
rect 227720 198500 227772 198552
rect 234528 198500 234580 198552
rect 267372 198500 267424 198552
rect 269028 198500 269080 198552
rect 282276 198500 282328 198552
rect 298376 198500 298428 198552
rect 302516 198500 302568 198552
rect 311808 198500 311860 198552
rect 330484 198500 330536 198552
rect 332968 198500 333020 198552
rect 340236 198500 340288 198552
rect 350448 198500 350500 198552
rect 420368 198500 420420 198552
rect 420828 198500 420880 198552
rect 58624 198432 58676 198484
rect 184204 198432 184256 198484
rect 184296 198432 184348 198484
rect 193588 198432 193640 198484
rect 195244 198432 195296 198484
rect 51724 198364 51776 198416
rect 181076 198364 181128 198416
rect 185584 198364 185636 198416
rect 196532 198364 196584 198416
rect 57244 198296 57296 198348
rect 189080 198296 189132 198348
rect 193864 198296 193916 198348
rect 214012 198432 214064 198484
rect 214656 198432 214708 198484
rect 226524 198432 226576 198484
rect 231768 198432 231820 198484
rect 266360 198432 266412 198484
rect 270408 198432 270460 198484
rect 283380 198432 283432 198484
rect 320088 198432 320140 198484
rect 338764 198432 338816 198484
rect 353760 198432 353812 198484
rect 429200 198432 429252 198484
rect 216772 198364 216824 198416
rect 227628 198364 227680 198416
rect 264980 198364 265032 198416
rect 267648 198364 267700 198416
rect 281724 198364 281776 198416
rect 299296 198364 299348 198416
rect 305184 198364 305236 198416
rect 344376 198364 344428 198416
rect 352564 198364 352616 198416
rect 356888 198364 356940 198416
rect 436100 198364 436152 198416
rect 196808 198296 196860 198348
rect 218244 198296 218296 198348
rect 223488 198296 223540 198348
rect 262772 198296 262824 198348
rect 268936 198296 268988 198348
rect 282920 198296 282972 198348
rect 326896 198296 326948 198348
rect 353944 198296 353996 198348
rect 35164 198228 35216 198280
rect 178040 198228 178092 198280
rect 178684 198228 178736 198280
rect 219440 198228 219492 198280
rect 220728 198228 220780 198280
rect 261668 198228 261720 198280
rect 264888 198228 264940 198280
rect 280804 198228 280856 198280
rect 285588 198228 285640 198280
rect 290096 198228 290148 198280
rect 315948 198228 316000 198280
rect 327908 198228 327960 198280
rect 330944 198228 330996 198280
rect 355784 198228 355836 198280
rect 358176 198228 358228 198280
rect 359832 198296 359884 198348
rect 443000 198296 443052 198348
rect 361028 198228 361080 198280
rect 362868 198228 362920 198280
rect 449900 198228 449952 198280
rect 29644 198160 29696 198212
rect 173992 198160 174044 198212
rect 184388 198160 184440 198212
rect 216220 198160 216272 198212
rect 217968 198160 218020 198212
rect 260196 198160 260248 198212
rect 262956 198160 263008 198212
rect 279700 198160 279752 198212
rect 304080 198160 304132 198212
rect 312544 198160 312596 198212
rect 318524 198160 318576 198212
rect 349344 198160 349396 198212
rect 351828 198160 351880 198212
rect 359464 198160 359516 198212
rect 18604 198092 18656 198144
rect 170220 198092 170272 198144
rect 191104 198092 191156 198144
rect 207388 198092 207440 198144
rect 213828 198092 213880 198144
rect 258540 198092 258592 198144
rect 260656 198092 260708 198144
rect 278780 198092 278832 198144
rect 285496 198092 285548 198144
rect 289820 198092 289872 198144
rect 309784 198092 309836 198144
rect 310428 198092 310480 198144
rect 11704 198024 11756 198076
rect 167644 198024 167696 198076
rect 184204 198024 184256 198076
rect 190460 198024 190512 198076
rect 192484 198024 192536 198076
rect 210516 198024 210568 198076
rect 210976 198024 211028 198076
rect 257068 198024 257120 198076
rect 259368 198024 259420 198076
rect 278228 198024 278280 198076
rect 278688 198024 278740 198076
rect 287060 198024 287112 198076
rect 302608 198024 302660 198076
rect 311992 198024 312044 198076
rect 323124 198092 323176 198144
rect 327448 198092 327500 198144
rect 358820 198092 358872 198144
rect 14464 197956 14516 198008
rect 169760 197956 169812 198008
rect 170404 197956 170456 198008
rect 180800 197956 180852 198008
rect 182824 197956 182876 198008
rect 187332 197956 187384 198008
rect 189724 197956 189776 198008
rect 204260 197956 204312 198008
rect 206928 197956 206980 198008
rect 255412 197956 255464 198008
rect 255964 197956 256016 198008
rect 275652 197956 275704 198008
rect 276664 197956 276716 198008
rect 285680 197956 285732 198008
rect 286968 197956 287020 198008
rect 290556 197956 290608 198008
rect 295800 197956 295852 198008
rect 296628 197956 296680 198008
rect 307208 197956 307260 198008
rect 317328 198024 317380 198076
rect 318064 198024 318116 198076
rect 357808 198024 357860 198076
rect 314016 197956 314068 198008
rect 314568 197956 314620 198008
rect 94504 197888 94556 197940
rect 205916 197888 205968 197940
rect 209044 197888 209096 197940
rect 241060 197888 241112 197940
rect 241428 197888 241480 197940
rect 270592 197888 270644 197940
rect 310336 197888 310388 197940
rect 327724 197956 327776 198008
rect 329748 197956 329800 198008
rect 363696 198092 363748 198144
rect 366916 198160 366968 198212
rect 385592 198160 385644 198212
rect 392400 198160 392452 198212
rect 482376 198160 482428 198212
rect 370596 198092 370648 198144
rect 366088 198024 366140 198076
rect 456800 198092 456852 198144
rect 370872 198024 370924 198076
rect 467840 198024 467892 198076
rect 360936 197956 360988 198008
rect 371976 197956 372028 198008
rect 373816 197956 373868 198008
rect 474740 197956 474792 198008
rect 339224 197888 339276 197940
rect 367744 197888 367796 197940
rect 369216 197888 369268 197940
rect 393964 197888 394016 197940
rect 101588 197820 101640 197872
rect 208952 197820 209004 197872
rect 209136 197820 209188 197872
rect 239404 197820 239456 197872
rect 253848 197820 253900 197872
rect 276204 197820 276256 197872
rect 298008 197820 298060 197872
rect 298744 197820 298796 197872
rect 322112 197820 322164 197872
rect 322848 197820 322900 197872
rect 328920 197820 328972 197872
rect 329748 197820 329800 197872
rect 333520 197820 333572 197872
rect 360936 197820 360988 197872
rect 367560 197820 367612 197872
rect 107568 197752 107620 197804
rect 212172 197752 212224 197804
rect 214564 197752 214616 197804
rect 225052 197752 225104 197804
rect 232504 197752 232556 197804
rect 261116 197752 261168 197804
rect 268384 197752 268436 197804
rect 277676 197752 277728 197804
rect 326344 197752 326396 197804
rect 340144 197752 340196 197804
rect 342168 197752 342220 197804
rect 367836 197752 367888 197804
rect 370136 197820 370188 197872
rect 394976 197820 395028 197872
rect 395896 197820 395948 197872
rect 378784 197752 378836 197804
rect 403624 197888 403676 197940
rect 467104 197888 467156 197940
rect 397000 197820 397052 197872
rect 114468 197684 114520 197736
rect 215300 197684 215352 197736
rect 216036 197684 216088 197736
rect 236276 197684 236328 197736
rect 251824 197684 251876 197736
rect 272524 197684 272576 197736
rect 306656 197684 306708 197736
rect 307668 197684 307720 197736
rect 310888 197684 310940 197736
rect 311808 197684 311860 197736
rect 320640 197684 320692 197736
rect 321468 197684 321520 197736
rect 328276 197684 328328 197736
rect 341524 197684 341576 197736
rect 343272 197684 343324 197736
rect 343456 197684 343508 197736
rect 348976 197684 349028 197736
rect 358084 197684 358136 197736
rect 359372 197684 359424 197736
rect 371884 197684 371936 197736
rect 376668 197684 376720 197736
rect 400864 197752 400916 197804
rect 403256 197820 403308 197872
rect 472624 197820 472676 197872
rect 409512 197752 409564 197804
rect 478144 197752 478196 197804
rect 380072 197684 380124 197736
rect 98644 197616 98696 197668
rect 198188 197616 198240 197668
rect 199384 197616 199436 197668
rect 211620 197616 211672 197668
rect 213184 197616 213236 197668
rect 236000 197616 236052 197668
rect 246304 197616 246356 197668
rect 259644 197616 259696 197668
rect 260748 197616 260800 197668
rect 279148 197616 279200 197668
rect 358360 197616 358412 197668
rect 364892 197616 364944 197668
rect 365536 197616 365588 197668
rect 372068 197616 372120 197668
rect 372344 197616 372396 197668
rect 381452 197616 381504 197668
rect 383200 197616 383252 197668
rect 405464 197684 405516 197736
rect 405648 197684 405700 197736
rect 412548 197684 412600 197736
rect 479524 197684 479576 197736
rect 105544 197548 105596 197600
rect 201500 197548 201552 197600
rect 215944 197548 215996 197600
rect 222200 197548 222252 197600
rect 224224 197548 224276 197600
rect 243084 197548 243136 197600
rect 125508 197480 125560 197532
rect 219900 197480 219952 197532
rect 256056 197480 256108 197532
rect 263140 197548 263192 197600
rect 267096 197548 267148 197600
rect 271420 197548 271472 197600
rect 300768 197548 300820 197600
rect 305644 197548 305696 197600
rect 309048 197548 309100 197600
rect 309876 197548 309928 197600
rect 312360 197548 312412 197600
rect 313924 197548 313976 197600
rect 321100 197548 321152 197600
rect 321376 197548 321428 197600
rect 325424 197548 325476 197600
rect 325608 197548 325660 197600
rect 364156 197548 364208 197600
rect 376024 197548 376076 197600
rect 384672 197548 384724 197600
rect 388444 197548 388496 197600
rect 260104 197480 260156 197532
rect 111064 197412 111116 197464
rect 173164 197344 173216 197396
rect 177580 197344 177632 197396
rect 181444 197344 181496 197396
rect 185308 197344 185360 197396
rect 186964 197344 187016 197396
rect 199660 197344 199712 197396
rect 202144 197412 202196 197464
rect 208492 197412 208544 197464
rect 264244 197412 264296 197464
rect 265716 197412 265768 197464
rect 269948 197480 270000 197532
rect 296352 197480 296404 197532
rect 298100 197480 298152 197532
rect 302056 197480 302108 197532
rect 304264 197480 304316 197532
rect 315488 197480 315540 197532
rect 318156 197480 318208 197532
rect 324228 197480 324280 197532
rect 356704 197480 356756 197532
rect 358820 197480 358872 197532
rect 359556 197480 359608 197532
rect 362408 197480 362460 197532
rect 366364 197480 366416 197532
rect 371792 197480 371844 197532
rect 385684 197480 385736 197532
rect 386144 197480 386196 197532
rect 389088 197480 389140 197532
rect 396724 197548 396776 197600
rect 399208 197548 399260 197600
rect 400128 197548 400180 197600
rect 406476 197616 406528 197668
rect 406568 197616 406620 197668
rect 407764 197548 407816 197600
rect 407856 197548 407908 197600
rect 409144 197548 409196 197600
rect 410892 197548 410944 197600
rect 411168 197548 411220 197600
rect 415308 197616 415360 197668
rect 269764 197412 269816 197464
rect 271972 197412 272024 197464
rect 282184 197412 282236 197464
rect 284852 197412 284904 197464
rect 284944 197412 284996 197464
rect 286508 197412 286560 197464
rect 300032 197412 300084 197464
rect 300768 197412 300820 197464
rect 301504 197412 301556 197464
rect 307024 197412 307076 197464
rect 314936 197412 314988 197464
rect 316684 197412 316736 197464
rect 323216 197412 323268 197464
rect 324136 197412 324188 197464
rect 332048 197412 332100 197464
rect 332508 197412 332560 197464
rect 334624 197412 334676 197464
rect 335176 197412 335228 197464
rect 336096 197412 336148 197464
rect 341616 197412 341668 197464
rect 345480 197412 345532 197464
rect 346216 197412 346268 197464
rect 351184 197412 351236 197464
rect 356796 197412 356848 197464
rect 361488 197412 361540 197464
rect 363604 197412 363656 197464
rect 364064 197412 364116 197464
rect 370688 197412 370740 197464
rect 373264 197412 373316 197464
rect 374644 197412 374696 197464
rect 374920 197412 374972 197464
rect 377404 197412 377456 197464
rect 387708 197412 387760 197464
rect 388536 197412 388588 197464
rect 389824 197412 389876 197464
rect 390468 197412 390520 197464
rect 398656 197480 398708 197532
rect 399484 197480 399536 197532
rect 402152 197480 402204 197532
rect 402888 197480 402940 197532
rect 403808 197480 403860 197532
rect 404268 197480 404320 197532
rect 404912 197480 404964 197532
rect 406384 197480 406436 197532
rect 407488 197480 407540 197532
rect 408316 197480 408368 197532
rect 408960 197480 409012 197532
rect 409696 197480 409748 197532
rect 410432 197480 410484 197532
rect 410984 197480 411036 197532
rect 412088 197480 412140 197532
rect 412548 197480 412600 197532
rect 418896 197480 418948 197532
rect 422300 197480 422352 197532
rect 202972 197344 203024 197396
rect 204904 197344 204956 197396
rect 205640 197344 205692 197396
rect 206284 197344 206336 197396
rect 207020 197344 207072 197396
rect 220176 197344 220228 197396
rect 223948 197344 224000 197396
rect 244924 197344 244976 197396
rect 247684 197344 247736 197396
rect 250444 197344 250496 197396
rect 253940 197344 253992 197396
rect 262864 197344 262916 197396
rect 264336 197344 264388 197396
rect 267004 197344 267056 197396
rect 269120 197344 269172 197396
rect 269856 197344 269908 197396
rect 270868 197344 270920 197396
rect 271144 197344 271196 197396
rect 273628 197344 273680 197396
rect 273904 197344 273956 197396
rect 275100 197344 275152 197396
rect 280804 197344 280856 197396
rect 281540 197344 281592 197396
rect 282276 197344 282328 197396
rect 284300 197344 284352 197396
rect 286324 197344 286376 197396
rect 287428 197344 287480 197396
rect 287704 197344 287756 197396
rect 289084 197344 289136 197396
rect 289728 197344 289780 197396
rect 291660 197344 291712 197396
rect 297456 197344 297508 197396
rect 298836 197344 298888 197396
rect 298928 197344 298980 197396
rect 300124 197344 300176 197396
rect 305736 197344 305788 197396
rect 306196 197344 306248 197396
rect 308312 197344 308364 197396
rect 309784 197344 309836 197396
rect 316592 197344 316644 197396
rect 317328 197344 317380 197396
rect 317972 197344 318024 197396
rect 318708 197344 318760 197396
rect 319536 197344 319588 197396
rect 322204 197344 322256 197396
rect 323768 197344 323820 197396
rect 324228 197344 324280 197396
rect 324872 197344 324924 197396
rect 325424 197344 325476 197396
rect 327816 197344 327868 197396
rect 328368 197344 328420 197396
rect 330392 197344 330444 197396
rect 331128 197344 331180 197396
rect 331496 197344 331548 197396
rect 332324 197344 332376 197396
rect 334992 197344 335044 197396
rect 335268 197344 335320 197396
rect 337200 197344 337252 197396
rect 338028 197344 338080 197396
rect 338672 197344 338724 197396
rect 339316 197344 339368 197396
rect 341248 197344 341300 197396
rect 342168 197344 342220 197396
rect 342904 197344 342956 197396
rect 343548 197344 343600 197396
rect 346032 197344 346084 197396
rect 346308 197344 346360 197396
rect 346952 197344 347004 197396
rect 347596 197344 347648 197396
rect 348608 197344 348660 197396
rect 349068 197344 349120 197396
rect 349528 197344 349580 197396
rect 350356 197344 350408 197396
rect 352656 197344 352708 197396
rect 353116 197344 353168 197396
rect 355232 197344 355284 197396
rect 360844 197344 360896 197396
rect 362040 197344 362092 197396
rect 362868 197344 362920 197396
rect 363512 197344 363564 197396
rect 364248 197344 364300 197396
rect 364984 197344 365036 197396
rect 365628 197344 365680 197396
rect 368388 197344 368440 197396
rect 370504 197344 370556 197396
rect 374368 197344 374420 197396
rect 375196 197344 375248 197396
rect 375840 197344 375892 197396
rect 376392 197344 376444 197396
rect 377496 197344 377548 197396
rect 377956 197344 378008 197396
rect 378416 197344 378468 197396
rect 379244 197344 379296 197396
rect 381544 197344 381596 197396
rect 382096 197344 382148 197396
rect 382648 197344 382700 197396
rect 383568 197344 383620 197396
rect 384120 197344 384172 197396
rect 384948 197344 385000 197396
rect 385776 197344 385828 197396
rect 386328 197344 386380 197396
rect 388352 197344 388404 197396
rect 388812 197344 388864 197396
rect 390928 197344 390980 197396
rect 392584 197344 392636 197396
rect 393044 197344 393096 197396
rect 393228 197344 393280 197396
rect 394056 197344 394108 197396
rect 395344 197344 395396 197396
rect 396632 197344 396684 197396
rect 397276 197344 397328 197396
rect 398104 197344 398156 197396
rect 398748 197344 398800 197396
rect 399576 197344 399628 197396
rect 400036 197344 400088 197396
rect 400680 197344 400732 197396
rect 401416 197344 401468 197396
rect 413008 197344 413060 197396
rect 413836 197344 413888 197396
rect 414664 197344 414716 197396
rect 415308 197344 415360 197396
rect 416136 197344 416188 197396
rect 416688 197344 416740 197396
rect 417240 197412 417292 197464
rect 418804 197412 418856 197464
rect 474004 197548 474056 197600
rect 482284 197480 482336 197532
rect 417424 197344 417476 197396
rect 417792 197344 417844 197396
rect 418068 197344 418120 197396
rect 418712 197344 418764 197396
rect 486424 197344 486476 197396
rect 200764 196868 200816 196920
rect 242992 196868 243044 196920
rect 169576 196800 169628 196852
rect 238944 196800 238996 196852
rect 88248 196732 88300 196784
rect 203892 196732 203944 196784
rect 380624 196732 380676 196784
rect 489920 196732 489972 196784
rect 39304 196664 39356 196716
rect 182180 196664 182232 196716
rect 188344 196664 188396 196716
rect 247132 196664 247184 196716
rect 386696 196664 386748 196716
rect 505100 196664 505152 196716
rect 14556 196596 14608 196648
rect 171324 196596 171376 196648
rect 180064 196596 180116 196648
rect 243636 196596 243688 196648
rect 391848 196596 391900 196648
rect 516140 196596 516192 196648
rect 165620 195236 165672 195288
rect 166172 195236 166224 195288
rect 172704 195236 172756 195288
rect 173348 195236 173400 195288
rect 178132 195236 178184 195288
rect 179052 195236 179104 195288
rect 182272 195236 182324 195288
rect 183100 195236 183152 195288
rect 186412 195236 186464 195288
rect 186780 195236 186832 195288
rect 237380 195236 237432 195288
rect 237932 195236 237984 195288
rect 251272 195236 251324 195288
rect 251916 195236 251968 195288
rect 254032 195236 254084 195288
rect 254860 195236 254912 195288
rect 190552 195032 190604 195084
rect 191380 195032 191432 195084
rect 245752 194488 245804 194540
rect 246212 194488 246264 194540
rect 244280 193264 244332 193316
rect 244648 193264 244700 193316
rect 428648 193128 428700 193180
rect 580172 193128 580224 193180
rect 168380 191972 168432 192024
rect 169300 191972 169352 192024
rect 198924 191224 198976 191276
rect 231860 191088 231912 191140
rect 232780 191088 232832 191140
rect 198924 191020 198976 191072
rect 244372 190884 244424 190936
rect 245108 190884 245160 190936
rect 2780 188844 2832 188896
rect 4804 188844 4856 188896
rect 198832 188368 198884 188420
rect 199016 188368 199068 188420
rect 209688 177284 209740 177336
rect 256792 177284 256844 177336
rect 258724 176672 258776 176724
rect 266544 176672 266596 176724
rect 220084 171776 220136 171828
rect 258172 171776 258224 171828
rect 424416 166948 424468 167000
rect 580172 166948 580224 167000
rect 3332 164160 3384 164212
rect 10416 164160 10468 164212
rect 204996 155184 205048 155236
rect 244464 155184 244516 155236
rect 428556 153144 428608 153196
rect 580172 153144 580224 153196
rect 3608 150356 3660 150408
rect 100116 150356 100168 150408
rect 429844 139340 429896 139392
rect 580172 139340 580224 139392
rect 421840 126896 421892 126948
rect 580172 126896 580224 126948
rect 425796 113092 425848 113144
rect 579804 113092 579856 113144
rect 3516 110712 3568 110764
rect 7656 110712 7708 110764
rect 428464 100648 428516 100700
rect 580172 100648 580224 100700
rect 3516 97928 3568 97980
rect 101496 97928 101548 97980
rect 103428 89156 103480 89208
rect 210056 89156 210108 89208
rect 81348 89088 81400 89140
rect 200212 89088 200264 89140
rect 35808 89020 35860 89072
rect 170404 89020 170456 89072
rect 23388 88952 23440 89004
rect 175464 88952 175516 89004
rect 384856 88952 384908 89004
rect 500960 88952 501012 89004
rect 135168 87728 135220 87780
rect 220176 87728 220228 87780
rect 43444 87660 43496 87712
rect 183652 87660 183704 87712
rect 28908 87592 28960 87644
rect 173164 87592 173216 87644
rect 242164 87592 242216 87644
rect 265164 87592 265216 87644
rect 372068 87592 372120 87644
rect 456892 87592 456944 87644
rect 421748 86912 421800 86964
rect 580172 86912 580224 86964
rect 341616 86504 341668 86556
rect 389180 86504 389232 86556
rect 366364 86436 366416 86488
rect 448520 86436 448572 86488
rect 362868 86368 362920 86420
rect 448612 86368 448664 86420
rect 379244 86300 379296 86352
rect 485780 86300 485832 86352
rect 106188 86232 106240 86284
rect 199384 86232 199436 86284
rect 206376 86232 206428 86284
rect 252744 86232 252796 86284
rect 340236 86232 340288 86284
rect 382372 86232 382424 86284
rect 388536 86232 388588 86284
rect 506480 86232 506532 86284
rect 3516 85484 3568 85536
rect 64144 85484 64196 85536
rect 162768 85076 162820 85128
rect 216036 85076 216088 85128
rect 143448 85008 143500 85060
rect 217324 85008 217376 85060
rect 113088 84940 113140 84992
rect 198004 84940 198056 84992
rect 198096 84940 198148 84992
rect 251364 84940 251416 84992
rect 137928 84872 137980 84924
rect 225052 84872 225104 84924
rect 370688 84872 370740 84924
rect 452660 84872 452712 84924
rect 95148 84804 95200 84856
rect 206284 84804 206336 84856
rect 400864 84804 400916 84856
rect 503720 84804 503772 84856
rect 147588 80656 147640 80708
rect 213276 80656 213328 80708
rect 424324 73108 424376 73160
rect 580172 73108 580224 73160
rect 3516 71612 3568 71664
rect 7564 71612 7616 71664
rect 425704 60664 425756 60716
rect 580172 60664 580224 60716
rect 3056 59304 3108 59356
rect 100024 59304 100076 59356
rect 421656 46860 421708 46912
rect 580172 46860 580224 46912
rect 3516 45500 3568 45552
rect 82084 45500 82136 45552
rect 99288 44820 99340 44872
rect 202144 44820 202196 44872
rect 385776 44820 385828 44872
rect 470600 44820 470652 44872
rect 370596 35164 370648 35216
rect 438860 35164 438912 35216
rect 2872 33056 2924 33108
rect 10324 33056 10376 33108
rect 508504 33056 508556 33108
rect 580172 33056 580224 33108
rect 388444 26868 388496 26920
rect 499580 26868 499632 26920
rect 370504 25508 370556 25560
rect 463700 25508 463752 25560
rect 392584 24080 392636 24132
rect 514760 24080 514812 24132
rect 245016 22856 245068 22908
rect 267832 22856 267884 22908
rect 216588 22788 216640 22840
rect 246304 22788 246356 22840
rect 32404 22720 32456 22772
rect 178132 22720 178184 22772
rect 202788 22720 202840 22772
rect 250444 22720 250496 22772
rect 395344 22720 395396 22772
rect 521660 22720 521712 22772
rect 382096 21360 382148 21412
rect 492680 21360 492732 21412
rect 3516 20612 3568 20664
rect 101404 20612 101456 20664
rect 421564 20612 421616 20664
rect 579988 20612 580040 20664
rect 356796 19932 356848 19984
rect 423680 19932 423732 19984
rect 140688 18572 140740 18624
rect 214656 18572 214708 18624
rect 161388 17484 161440 17536
rect 213184 17484 213236 17536
rect 144828 17416 144880 17468
rect 227812 17416 227864 17468
rect 129648 17348 129700 17400
rect 215944 17348 215996 17400
rect 110328 17280 110380 17332
rect 196716 17280 196768 17332
rect 196808 17280 196860 17332
rect 244372 17280 244424 17332
rect 354496 17280 354548 17332
rect 430580 17280 430632 17332
rect 133788 17212 133840 17264
rect 223672 17212 223724 17264
rect 341524 17212 341576 17264
rect 371240 17212 371292 17264
rect 407764 17212 407816 17264
rect 496820 17212 496872 17264
rect 124128 16192 124180 16244
rect 178684 16192 178736 16244
rect 396724 16192 396776 16244
rect 467104 16192 467156 16244
rect 119896 16124 119948 16176
rect 177304 16124 177356 16176
rect 371884 16124 371936 16176
rect 442632 16124 442684 16176
rect 165528 16056 165580 16108
rect 237472 16056 237524 16108
rect 371976 16056 372028 16108
rect 445760 16056 445812 16108
rect 139308 15988 139360 16040
rect 226432 15988 226484 16040
rect 377956 15988 378008 16040
rect 484032 15988 484084 16040
rect 92388 15920 92440 15972
rect 204904 15920 204956 15972
rect 417424 15920 417476 15972
rect 525432 15920 525484 15972
rect 45468 15852 45520 15904
rect 181444 15852 181496 15904
rect 205088 15852 205140 15904
rect 248696 15852 248748 15904
rect 388996 15852 389048 15904
rect 508872 15852 508924 15904
rect 357348 14764 357400 14816
rect 437480 14764 437532 14816
rect 117228 14696 117280 14748
rect 184388 14696 184440 14748
rect 406476 14696 406528 14748
rect 490012 14696 490064 14748
rect 166908 14628 166960 14680
rect 237380 14628 237432 14680
rect 318156 14628 318208 14680
rect 341984 14628 342036 14680
rect 418896 14628 418948 14680
rect 511264 14628 511316 14680
rect 126888 14560 126940 14612
rect 219716 14560 219768 14612
rect 324136 14560 324188 14612
rect 358268 14560 358320 14612
rect 390376 14560 390428 14612
rect 513564 14560 513616 14612
rect 85488 14492 85540 14544
rect 201776 14492 201828 14544
rect 238024 14492 238076 14544
rect 263692 14492 263744 14544
rect 321284 14492 321336 14544
rect 356336 14492 356388 14544
rect 361028 14492 361080 14544
rect 377680 14492 377732 14544
rect 395896 14492 395948 14544
rect 522304 14492 522356 14544
rect 19248 14424 19300 14476
rect 172704 14424 172756 14476
rect 202144 14424 202196 14476
rect 245752 14424 245804 14476
rect 246948 14424 247000 14476
rect 273352 14424 273404 14476
rect 329656 14424 329708 14476
rect 367928 14424 367980 14476
rect 393136 14424 393188 14476
rect 520280 14424 520332 14476
rect 145932 13132 145984 13184
rect 229192 13132 229244 13184
rect 131028 13064 131080 13116
rect 222292 13064 222344 13116
rect 251088 13064 251140 13116
rect 274824 13064 274876 13116
rect 358728 13064 358780 13116
rect 441528 13064 441580 13116
rect 325424 11840 325476 11892
rect 363512 11772 363564 11824
rect 379336 11772 379388 11824
rect 487160 11772 487212 11824
rect 328368 11704 328420 11756
rect 370136 11704 370188 11756
rect 382188 11704 382240 11756
rect 494704 11704 494756 11756
rect 358176 10412 358228 10464
rect 433984 10412 434036 10464
rect 367836 10344 367888 10396
rect 403624 10344 403676 10396
rect 403716 10344 403768 10396
rect 482100 10344 482152 10396
rect 363696 10276 363748 10328
rect 375104 10276 375156 10328
rect 374644 10208 374696 10260
rect 473912 10276 473964 10328
rect 175464 9528 175516 9580
rect 241612 9528 241664 9580
rect 171968 9460 172020 9512
rect 240232 9460 240284 9512
rect 136456 9392 136508 9444
rect 214564 9392 214616 9444
rect 135260 9324 135312 9376
rect 223856 9324 223908 9376
rect 350356 9324 350408 9376
rect 420184 9324 420236 9376
rect 131764 9256 131816 9308
rect 222384 9256 222436 9308
rect 353116 9256 353168 9308
rect 427268 9256 427320 9308
rect 77392 9188 77444 9240
rect 198832 9188 198884 9240
rect 385684 9188 385736 9240
rect 460388 9188 460440 9240
rect 73804 9120 73856 9172
rect 197636 9120 197688 9172
rect 360108 9120 360160 9172
rect 445024 9120 445076 9172
rect 70308 9052 70360 9104
rect 196072 9052 196124 9104
rect 377404 9052 377456 9104
rect 478052 9052 478104 9104
rect 66720 8984 66772 9036
rect 194692 8984 194744 9036
rect 376576 8984 376628 9036
rect 480536 8984 480588 9036
rect 482376 8984 482428 9036
rect 518348 8984 518400 9036
rect 63224 8916 63276 8968
rect 193312 8916 193364 8968
rect 383476 8916 383528 8968
rect 498200 8916 498252 8968
rect 108120 8236 108172 8288
rect 212632 8236 212684 8288
rect 401324 8236 401376 8288
rect 538404 8236 538456 8288
rect 104532 8168 104584 8220
rect 211344 8168 211396 8220
rect 402796 8168 402848 8220
rect 541992 8168 542044 8220
rect 101036 8100 101088 8152
rect 209964 8100 210016 8152
rect 404176 8100 404228 8152
rect 545488 8100 545540 8152
rect 97448 8032 97500 8084
rect 207204 8032 207256 8084
rect 405556 8032 405608 8084
rect 549076 8032 549128 8084
rect 93952 7964 94004 8016
rect 205824 7964 205876 8016
rect 408316 7964 408368 8016
rect 552664 7964 552716 8016
rect 90364 7896 90416 7948
rect 204352 7896 204404 7948
rect 409696 7896 409748 7948
rect 556160 7896 556212 7948
rect 86868 7828 86920 7880
rect 203064 7828 203116 7880
rect 410984 7828 411036 7880
rect 559748 7828 559800 7880
rect 59636 7760 59688 7812
rect 190552 7760 190604 7812
rect 412548 7760 412600 7812
rect 563244 7760 563296 7812
rect 56048 7692 56100 7744
rect 189356 7692 189408 7744
rect 413744 7692 413796 7744
rect 566832 7692 566884 7744
rect 52552 7624 52604 7676
rect 187792 7624 187844 7676
rect 415216 7624 415268 7676
rect 570328 7624 570380 7676
rect 48964 7556 49016 7608
rect 186412 7556 186464 7608
rect 416596 7556 416648 7608
rect 573916 7556 573968 7608
rect 111616 7488 111668 7540
rect 214104 7488 214156 7540
rect 400036 7488 400088 7540
rect 534908 7488 534960 7540
rect 115204 7420 115256 7472
rect 215576 7420 215628 7472
rect 398748 7420 398800 7472
rect 531320 7420 531372 7472
rect 118792 7352 118844 7404
rect 216772 7352 216824 7404
rect 397276 7352 397328 7404
rect 527824 7352 527876 7404
rect 122288 7284 122340 7336
rect 218244 7284 218296 7336
rect 355968 7284 356020 7336
rect 435548 7284 435600 7336
rect 149520 7216 149572 7268
rect 230664 7216 230716 7268
rect 354588 7216 354640 7268
rect 432052 7216 432104 7268
rect 153016 7148 153068 7200
rect 232136 7148 232188 7200
rect 353208 7148 353260 7200
rect 428464 7148 428516 7200
rect 156604 7080 156656 7132
rect 233332 7080 233384 7132
rect 351828 7080 351880 7132
rect 424968 7080 425020 7132
rect 160100 7012 160152 7064
rect 234804 7012 234856 7064
rect 350448 7012 350500 7064
rect 421380 7012 421432 7064
rect 83280 6808 83332 6860
rect 201684 6808 201736 6860
rect 447784 6808 447836 6860
rect 580172 6808 580224 6860
rect 79692 6740 79744 6792
rect 200120 6740 200172 6792
rect 376668 6740 376720 6792
rect 481732 6740 481784 6792
rect 44272 6672 44324 6724
rect 185032 6672 185084 6724
rect 378048 6672 378100 6724
rect 485228 6672 485280 6724
rect 40684 6604 40736 6656
rect 182272 6604 182324 6656
rect 205180 6604 205232 6656
rect 254032 6604 254084 6656
rect 379428 6604 379480 6656
rect 488816 6604 488868 6656
rect 37188 6536 37240 6588
rect 180984 6536 181036 6588
rect 201500 6536 201552 6588
rect 252836 6536 252888 6588
rect 380716 6536 380768 6588
rect 492312 6536 492364 6588
rect 33600 6468 33652 6520
rect 179512 6468 179564 6520
rect 197912 6468 197964 6520
rect 251272 6468 251324 6520
rect 383568 6468 383620 6520
rect 495900 6468 495952 6520
rect 30104 6400 30156 6452
rect 178224 6400 178276 6452
rect 194416 6400 194468 6452
rect 249892 6400 249944 6452
rect 384948 6400 385000 6452
rect 499396 6400 499448 6452
rect 26516 6332 26568 6384
rect 176936 6332 176988 6384
rect 190828 6332 190880 6384
rect 248512 6332 248564 6384
rect 386328 6332 386380 6384
rect 502984 6332 503036 6384
rect 21824 6264 21876 6316
rect 175372 6264 175424 6316
rect 187332 6264 187384 6316
rect 247224 6264 247276 6316
rect 338764 6264 338816 6316
rect 352840 6264 352892 6316
rect 387616 6264 387668 6316
rect 506480 6264 506532 6316
rect 8760 6196 8812 6248
rect 168380 6196 168432 6248
rect 170772 6196 170824 6248
rect 240324 6196 240376 6248
rect 340144 6196 340196 6248
rect 366916 6196 366968 6248
rect 389088 6196 389140 6248
rect 510068 6196 510120 6248
rect 4068 6128 4120 6180
rect 167092 6128 167144 6180
rect 167184 6128 167236 6180
rect 238760 6128 238812 6180
rect 317236 6128 317288 6180
rect 345756 6128 345808 6180
rect 367744 6128 367796 6180
rect 396540 6128 396592 6180
rect 417976 6128 418028 6180
rect 577412 6128 577464 6180
rect 128176 6060 128228 6112
rect 220912 6060 220964 6112
rect 372528 6060 372580 6112
rect 473452 6060 473504 6112
rect 141240 5992 141292 6044
rect 226524 5992 226576 6044
rect 375196 5992 375248 6044
rect 476948 5992 477000 6044
rect 144736 5924 144788 5976
rect 227996 5924 228048 5976
rect 371148 5924 371200 5976
rect 469864 5924 469916 5976
rect 148324 5856 148376 5908
rect 230572 5856 230624 5908
rect 369768 5856 369820 5908
rect 466276 5856 466328 5908
rect 151820 5788 151872 5840
rect 231952 5788 232004 5840
rect 368388 5788 368440 5840
rect 462780 5788 462832 5840
rect 155408 5720 155460 5772
rect 233240 5720 233292 5772
rect 367008 5720 367060 5772
rect 459192 5720 459244 5772
rect 158904 5652 158956 5704
rect 234712 5652 234764 5704
rect 365628 5652 365680 5704
rect 455696 5652 455748 5704
rect 163688 5584 163740 5636
rect 236276 5584 236328 5636
rect 364248 5584 364300 5636
rect 452108 5584 452160 5636
rect 62028 5448 62080 5500
rect 191932 5448 191984 5500
rect 221556 5448 221608 5500
rect 262404 5448 262456 5500
rect 339316 5448 339368 5500
rect 395344 5448 395396 5500
rect 402888 5448 402940 5500
rect 540796 5448 540848 5500
rect 58440 5380 58492 5432
rect 190644 5380 190696 5432
rect 218060 5380 218112 5432
rect 261024 5380 261076 5432
rect 340696 5380 340748 5432
rect 398932 5380 398984 5432
rect 404268 5380 404320 5432
rect 544384 5380 544436 5432
rect 54944 5312 54996 5364
rect 189264 5312 189316 5364
rect 214472 5312 214524 5364
rect 258264 5312 258316 5364
rect 340788 5312 340840 5364
rect 400128 5312 400180 5364
rect 405648 5312 405700 5364
rect 547880 5312 547932 5364
rect 51356 5244 51408 5296
rect 187700 5244 187752 5296
rect 211068 5244 211120 5296
rect 256884 5244 256936 5296
rect 307576 5244 307628 5296
rect 324412 5244 324464 5296
rect 342076 5244 342128 5296
rect 402520 5244 402572 5296
rect 407028 5244 407080 5296
rect 551468 5244 551520 5296
rect 47860 5176 47912 5228
rect 186504 5176 186556 5228
rect 207388 5176 207440 5228
rect 255412 5176 255464 5228
rect 309876 5176 309928 5228
rect 169668 5108 169720 5160
rect 209136 5108 209188 5160
rect 311808 5108 311860 5160
rect 327816 5176 327868 5228
rect 343272 5176 343324 5228
rect 343456 5176 343508 5228
rect 406016 5176 406068 5228
rect 408408 5176 408460 5228
rect 554964 5176 555016 5228
rect 12348 5040 12400 5092
rect 171232 5040 171284 5092
rect 173164 5040 173216 5092
rect 209044 5040 209096 5092
rect 313924 5040 313976 5092
rect 328000 5108 328052 5160
rect 344928 5108 344980 5160
rect 409604 5108 409656 5160
rect 409788 5108 409840 5160
rect 558552 5108 558604 5160
rect 331588 5040 331640 5092
rect 346216 5040 346268 5092
rect 410800 5040 410852 5092
rect 415308 5040 415360 5092
rect 7656 4972 7708 5024
rect 168472 4972 168524 5024
rect 196808 4972 196860 5024
rect 251456 4972 251508 5024
rect 311716 4972 311768 5024
rect 332692 4972 332744 5024
rect 343364 4972 343416 5024
rect 407212 4972 407264 5024
rect 411076 4972 411128 5024
rect 2872 4904 2924 4956
rect 167000 4904 167052 4956
rect 193220 4904 193272 4956
rect 249800 4904 249852 4956
rect 314568 4904 314620 4956
rect 338672 4904 338724 4956
rect 346124 4904 346176 4956
rect 413100 4904 413152 4956
rect 413836 4904 413888 4956
rect 416596 4904 416648 4956
rect 565636 5040 565688 5092
rect 562048 4972 562100 5024
rect 1676 4836 1728 4888
rect 165620 4836 165672 4888
rect 189724 4836 189776 4888
rect 248420 4836 248472 4888
rect 314476 4836 314528 4888
rect 339868 4836 339920 4888
rect 347688 4836 347740 4888
rect 416688 4836 416740 4888
rect 569132 4904 569184 4956
rect 572720 4836 572772 4888
rect 572 4768 624 4820
rect 165712 4768 165764 4820
rect 174268 4768 174320 4820
rect 241520 4768 241572 4820
rect 318064 4768 318116 4820
rect 346952 4768 347004 4820
rect 349068 4768 349120 4820
rect 417884 4768 417936 4820
rect 418068 4768 418120 4820
rect 576308 4768 576360 4820
rect 65524 4700 65576 4752
rect 193404 4700 193456 4752
rect 200304 4700 200356 4752
rect 252560 4700 252612 4752
rect 334992 4700 335044 4752
rect 337936 4700 337988 4752
rect 393044 4700 393096 4752
rect 401416 4700 401468 4752
rect 537208 4700 537260 4752
rect 72608 4632 72660 4684
rect 197544 4632 197596 4684
rect 203892 4632 203944 4684
rect 254124 4632 254176 4684
rect 335084 4632 335136 4684
rect 388260 4632 388312 4684
rect 400036 4632 400088 4684
rect 533712 4632 533764 4684
rect 69112 4564 69164 4616
rect 194784 4564 194836 4616
rect 338028 4564 338080 4616
rect 391848 4564 391900 4616
rect 397368 4564 397420 4616
rect 530124 4564 530176 4616
rect 76196 4496 76248 4548
rect 198924 4496 198976 4548
rect 335176 4496 335228 4548
rect 385960 4496 386012 4548
rect 395988 4496 396040 4548
rect 526628 4496 526680 4548
rect 126980 4428 127032 4480
rect 220820 4428 220872 4480
rect 333888 4428 333940 4480
rect 384764 4428 384816 4480
rect 394608 4428 394660 4480
rect 523040 4428 523092 4480
rect 150624 4360 150676 4412
rect 230756 4360 230808 4412
rect 332416 4360 332468 4412
rect 381176 4360 381228 4412
rect 393228 4360 393280 4412
rect 519544 4360 519596 4412
rect 154212 4292 154264 4344
rect 231860 4292 231912 4344
rect 332324 4292 332376 4344
rect 378876 4292 378928 4344
rect 391756 4292 391808 4344
rect 515956 4292 516008 4344
rect 157800 4224 157852 4276
rect 234620 4224 234672 4276
rect 367928 4224 367980 4276
rect 17040 4156 17092 4208
rect 172796 4156 172848 4208
rect 177856 4156 177908 4208
rect 224224 4156 224276 4208
rect 347596 4156 347648 4208
rect 11152 4020 11204 4072
rect 18604 4020 18656 4072
rect 20628 4020 20680 4072
rect 61384 4088 61436 4140
rect 64328 4088 64380 4140
rect 184296 4088 184348 4140
rect 242900 4088 242952 4140
rect 267096 4088 267148 4140
rect 281908 4088 281960 4140
rect 288532 4088 288584 4140
rect 296628 4088 296680 4140
rect 297272 4088 297324 4140
rect 303436 4088 303488 4140
rect 312544 4088 312596 4140
rect 316224 4088 316276 4140
rect 331128 4088 331180 4140
rect 390468 4224 390520 4276
rect 512460 4224 512512 4276
rect 414296 4156 414348 4208
rect 490748 4156 490800 4208
rect 374092 4088 374144 4140
rect 381544 4088 381596 4140
rect 472256 4088 472308 4140
rect 489920 4088 489972 4140
rect 491116 4088 491168 4140
rect 582196 4088 582248 4140
rect 35992 4020 36044 4072
rect 51724 4020 51776 4072
rect 53748 4020 53800 4072
rect 57152 4020 57204 4072
rect 57244 4020 57296 4072
rect 184204 4020 184256 4072
rect 228732 4020 228784 4072
rect 242164 4020 242216 4072
rect 244096 4020 244148 4072
rect 50160 3952 50212 4004
rect 46664 3884 46716 3936
rect 39580 3816 39632 3868
rect 185216 3952 185268 4004
rect 232228 3952 232280 4004
rect 267004 4020 267056 4072
rect 306196 4020 306248 4072
rect 319720 4020 319772 4072
rect 329748 4020 329800 4072
rect 372896 4020 372948 4072
rect 375288 4020 375340 4072
rect 479340 4020 479392 4072
rect 486424 4020 486476 4072
rect 578608 4020 578660 4072
rect 269764 3952 269816 4004
rect 306288 3952 306340 4004
rect 320916 3952 320968 4004
rect 332508 3952 332560 4004
rect 379980 3952 380032 4004
rect 399484 3952 399536 4004
rect 532516 3952 532568 4004
rect 192024 3884 192076 3936
rect 205088 3884 205140 3936
rect 225144 3884 225196 3936
rect 238024 3884 238076 3936
rect 241704 3884 241756 3936
rect 269856 3884 269908 3936
rect 300768 3884 300820 3936
rect 306748 3884 306800 3936
rect 313832 3884 313884 3936
rect 19432 3748 19484 3800
rect 29644 3748 29696 3800
rect 32496 3748 32548 3800
rect 182824 3816 182876 3868
rect 199108 3816 199160 3868
rect 206376 3816 206428 3868
rect 219256 3816 219308 3868
rect 232504 3816 232556 3868
rect 237012 3816 237064 3868
rect 67916 3680 67968 3732
rect 76564 3680 76616 3732
rect 80888 3680 80940 3732
rect 81348 3680 81400 3732
rect 84476 3680 84528 3732
rect 85488 3680 85540 3732
rect 91560 3680 91612 3732
rect 92388 3680 92440 3732
rect 92756 3680 92808 3732
rect 94504 3680 94556 3732
rect 98644 3680 98696 3732
rect 99288 3680 99340 3732
rect 99840 3680 99892 3732
rect 101588 3680 101640 3732
rect 102232 3680 102284 3732
rect 103428 3680 103480 3732
rect 105728 3680 105780 3732
rect 106188 3680 106240 3732
rect 106924 3680 106976 3732
rect 107568 3680 107620 3732
rect 109316 3680 109368 3732
rect 110328 3680 110380 3732
rect 114008 3680 114060 3732
rect 114468 3680 114520 3732
rect 116400 3680 116452 3732
rect 117228 3680 117280 3732
rect 123484 3680 123536 3732
rect 124128 3680 124180 3732
rect 124680 3680 124732 3732
rect 125508 3680 125560 3732
rect 125876 3680 125928 3732
rect 126888 3680 126940 3732
rect 130568 3680 130620 3732
rect 131028 3680 131080 3732
rect 132960 3680 133012 3732
rect 133788 3680 133840 3732
rect 134156 3680 134208 3732
rect 135168 3680 135220 3732
rect 138848 3680 138900 3732
rect 139308 3680 139360 3732
rect 140044 3680 140096 3732
rect 140688 3680 140740 3732
rect 142436 3680 142488 3732
rect 143448 3680 143500 3732
rect 143540 3680 143592 3732
rect 144828 3680 144880 3732
rect 147128 3680 147180 3732
rect 147588 3680 147640 3732
rect 168656 3680 168708 3732
rect 24216 3612 24268 3664
rect 175556 3612 175608 3664
rect 182364 3748 182416 3800
rect 184940 3748 184992 3800
rect 202144 3748 202196 3800
rect 223948 3748 224000 3800
rect 256056 3748 256108 3800
rect 264244 3816 264296 3868
rect 300676 3816 300728 3868
rect 307944 3816 307996 3868
rect 309784 3816 309836 3868
rect 325608 3884 325660 3936
rect 326804 3816 326856 3868
rect 176660 3680 176712 3732
rect 200764 3680 200816 3732
rect 229836 3680 229888 3732
rect 263048 3748 263100 3800
rect 280344 3748 280396 3800
rect 304908 3748 304960 3800
rect 318524 3748 318576 3800
rect 318708 3748 318760 3800
rect 179420 3612 179472 3664
rect 180248 3612 180300 3664
rect 204904 3612 204956 3664
rect 212172 3612 212224 3664
rect 220084 3612 220136 3664
rect 226340 3612 226392 3664
rect 262864 3680 262916 3732
rect 308956 3680 309008 3732
rect 258264 3612 258316 3664
rect 258724 3612 258776 3664
rect 265348 3612 265400 3664
rect 280804 3612 280856 3664
rect 284300 3612 284352 3664
rect 285496 3612 285548 3664
rect 305644 3612 305696 3664
rect 309048 3612 309100 3664
rect 313188 3680 313240 3732
rect 316684 3680 316736 3732
rect 329196 3816 329248 3868
rect 335268 3884 335320 3936
rect 387156 3884 387208 3936
rect 401508 3884 401560 3936
rect 539600 3884 539652 3936
rect 336648 3816 336700 3868
rect 390652 3816 390704 3868
rect 406384 3816 406436 3868
rect 546684 3816 546736 3868
rect 348056 3748 348108 3800
rect 352564 3748 352616 3800
rect 408408 3748 408460 3800
rect 409144 3748 409196 3800
rect 553768 3748 553820 3800
rect 327724 3680 327776 3732
rect 330392 3680 330444 3732
rect 330484 3680 330536 3732
rect 333888 3680 333940 3732
rect 342168 3680 342220 3732
rect 401324 3680 401376 3732
rect 411168 3680 411220 3732
rect 560852 3680 560904 3732
rect 337476 3612 337528 3664
rect 339408 3612 339460 3664
rect 397736 3612 397788 3664
rect 15936 3544 15988 3596
rect 172520 3544 172572 3596
rect 188528 3544 188580 3596
rect 244924 3544 244976 3596
rect 251180 3544 251232 3596
rect 273904 3544 273956 3596
rect 276020 3544 276072 3596
rect 277308 3544 277360 3596
rect 279516 3544 279568 3596
rect 286324 3544 286376 3596
rect 303528 3544 303580 3596
rect 5264 3476 5316 3528
rect 11704 3476 11756 3528
rect 13544 3476 13596 3528
rect 14556 3476 14608 3528
rect 14740 3476 14792 3528
rect 171324 3476 171376 3528
rect 179052 3476 179104 3528
rect 180064 3476 180116 3528
rect 6460 3408 6512 3460
rect 164884 3408 164936 3460
rect 165528 3408 165580 3460
rect 166080 3408 166132 3460
rect 166908 3408 166960 3460
rect 168380 3408 168432 3460
rect 169576 3408 169628 3460
rect 18236 3340 18288 3392
rect 19248 3340 19300 3392
rect 27712 3340 27764 3392
rect 28908 3340 28960 3392
rect 31300 3340 31352 3392
rect 32404 3340 32456 3392
rect 34796 3340 34848 3392
rect 35808 3340 35860 3392
rect 38384 3340 38436 3392
rect 39304 3340 39356 3392
rect 41880 3340 41932 3392
rect 43444 3340 43496 3392
rect 43076 3272 43128 3324
rect 58624 3340 58676 3392
rect 71504 3340 71556 3392
rect 185584 3476 185636 3528
rect 186136 3476 186188 3528
rect 188344 3476 188396 3528
rect 183744 3408 183796 3460
rect 240508 3476 240560 3528
rect 241428 3476 241480 3528
rect 246396 3476 246448 3528
rect 246948 3476 247000 3528
rect 247592 3476 247644 3528
rect 271144 3476 271196 3528
rect 271236 3476 271288 3528
rect 271788 3476 271840 3528
rect 274824 3476 274876 3528
rect 276664 3476 276716 3528
rect 277124 3476 277176 3528
rect 284944 3476 284996 3528
rect 288992 3476 289044 3528
rect 289728 3476 289780 3528
rect 291384 3476 291436 3528
rect 292488 3476 292540 3528
rect 294052 3476 294104 3528
rect 294880 3476 294932 3528
rect 300124 3476 300176 3528
rect 304356 3476 304408 3528
rect 307668 3544 307720 3596
rect 322112 3544 322164 3596
rect 322756 3544 322808 3596
rect 357716 3544 357768 3596
rect 358268 3544 358320 3596
rect 359924 3544 359976 3596
rect 418988 3544 419040 3596
rect 315028 3476 315080 3528
rect 317236 3476 317288 3528
rect 181444 3340 181496 3392
rect 244280 3408 244332 3460
rect 249984 3408 250036 3460
rect 251088 3408 251140 3460
rect 258172 3408 258224 3460
rect 258264 3408 258316 3460
rect 259368 3408 259420 3460
rect 259460 3408 259512 3460
rect 260564 3408 260616 3460
rect 261760 3408 261812 3460
rect 262956 3408 263008 3460
rect 264152 3408 264204 3460
rect 264888 3408 264940 3460
rect 266544 3408 266596 3460
rect 267648 3408 267700 3460
rect 273628 3408 273680 3460
rect 282184 3408 282236 3460
rect 296536 3408 296588 3460
rect 299664 3408 299716 3460
rect 304816 3408 304868 3460
rect 317328 3408 317380 3460
rect 340972 3476 341024 3528
rect 343548 3476 343600 3528
rect 404820 3476 404872 3528
rect 414664 3476 414716 3528
rect 415492 3476 415544 3528
rect 344560 3408 344612 3460
rect 346308 3408 346360 3460
rect 411904 3408 411956 3460
rect 413928 3408 413980 3460
rect 568028 3612 568080 3664
rect 419264 3544 419316 3596
rect 575112 3544 575164 3596
rect 420828 3476 420880 3528
rect 583392 3476 583444 3528
rect 419448 3408 419500 3460
rect 581000 3408 581052 3460
rect 206192 3340 206244 3392
rect 206928 3340 206980 3392
rect 208584 3340 208636 3392
rect 209688 3340 209740 3392
rect 209780 3340 209832 3392
rect 210976 3340 211028 3392
rect 213368 3340 213420 3392
rect 213828 3340 213880 3392
rect 215668 3340 215720 3392
rect 216588 3340 216640 3392
rect 216864 3340 216916 3392
rect 217968 3340 218020 3392
rect 222752 3340 222804 3392
rect 223488 3340 223540 3392
rect 231032 3340 231084 3392
rect 231768 3340 231820 3392
rect 233424 3340 233476 3392
rect 234528 3340 234580 3392
rect 235816 3340 235868 3392
rect 60832 3272 60884 3324
rect 71044 3272 71096 3324
rect 78588 3272 78640 3324
rect 186964 3272 187016 3324
rect 234620 3272 234672 3324
rect 235908 3272 235960 3324
rect 238116 3272 238168 3324
rect 238668 3272 238720 3324
rect 245844 3340 245896 3392
rect 254676 3340 254728 3392
rect 245016 3272 245068 3324
rect 245200 3272 245252 3324
rect 251824 3272 251876 3324
rect 255872 3272 255924 3324
rect 272432 3340 272484 3392
rect 282276 3340 282328 3392
rect 304264 3340 304316 3392
rect 311440 3340 311492 3392
rect 324228 3340 324280 3392
rect 361120 3340 361172 3392
rect 363604 3340 363656 3392
rect 447416 3340 447468 3392
rect 448520 3340 448572 3392
rect 449808 3340 449860 3392
rect 456800 3340 456852 3392
rect 458088 3340 458140 3392
rect 482192 3340 482244 3392
rect 571524 3340 571576 3392
rect 9956 3204 10008 3256
rect 14464 3204 14516 3256
rect 28908 3204 28960 3256
rect 35164 3204 35216 3256
rect 89168 3204 89220 3256
rect 189632 3204 189684 3256
rect 239312 3204 239364 3256
rect 260104 3204 260156 3256
rect 276204 3272 276256 3324
rect 280712 3272 280764 3324
rect 287336 3272 287388 3324
rect 310428 3272 310480 3324
rect 325424 3272 325476 3324
rect 365812 3272 365864 3324
rect 376484 3272 376536 3324
rect 378784 3272 378836 3324
rect 461584 3272 461636 3324
rect 479524 3272 479576 3324
rect 564440 3272 564492 3324
rect 277584 3204 277636 3256
rect 325516 3204 325568 3256
rect 364616 3204 364668 3256
rect 376024 3204 376076 3256
rect 454500 3204 454552 3256
rect 478236 3204 478288 3256
rect 557356 3204 557408 3256
rect 96252 3136 96304 3188
rect 191104 3136 191156 3188
rect 257068 3136 257120 3188
rect 268384 3136 268436 3188
rect 287796 3136 287848 3188
rect 291292 3136 291344 3188
rect 298744 3136 298796 3188
rect 301964 3136 302016 3188
rect 307024 3136 307076 3188
rect 310244 3136 310296 3188
rect 322848 3136 322900 3188
rect 357532 3136 357584 3188
rect 358176 3136 358228 3188
rect 360936 3136 360988 3188
rect 75000 3068 75052 3120
rect 98552 3068 98604 3120
rect 103336 3068 103388 3120
rect 192484 3068 192536 3120
rect 248788 3068 248840 3120
rect 273444 3068 273496 3120
rect 283104 3068 283156 3120
rect 287704 3068 287756 3120
rect 321376 3068 321428 3120
rect 355232 3068 355284 3120
rect 356704 3068 356756 3120
rect 362316 3068 362368 3120
rect 364984 3136 365036 3188
rect 440332 3136 440384 3188
rect 474004 3136 474056 3188
rect 550272 3136 550324 3188
rect 383568 3068 383620 3120
rect 393964 3068 394016 3120
rect 465172 3068 465224 3120
rect 472624 3068 472676 3120
rect 543188 3068 543240 3120
rect 82084 3000 82136 3052
rect 105544 3000 105596 3052
rect 110512 3000 110564 3052
rect 193864 3000 193916 3052
rect 252376 3000 252428 3052
rect 255964 3000 256016 3052
rect 298836 3000 298888 3052
rect 300768 3000 300820 3052
rect 321468 3000 321520 3052
rect 354036 3000 354088 3052
rect 360844 3000 360896 3052
rect 433248 3000 433300 3052
rect 471244 3000 471296 3052
rect 536104 3000 536156 3052
rect 85672 2932 85724 2984
rect 111064 2932 111116 2984
rect 117596 2932 117648 2984
rect 195244 2932 195296 2984
rect 195612 2932 195664 2984
rect 198096 2932 198148 2984
rect 290188 2932 290240 2984
rect 291476 2932 291528 2984
rect 322204 2932 322256 2984
rect 351644 2932 351696 2984
rect 359464 2932 359516 2984
rect 426164 2932 426216 2984
rect 467196 2932 467248 2984
rect 121092 2864 121144 2916
rect 196624 2864 196676 2916
rect 267740 2864 267792 2916
rect 269028 2864 269080 2916
rect 336004 2864 336056 2916
rect 350448 2864 350500 2916
rect 353944 2864 353996 2916
rect 368204 2864 368256 2916
rect 522304 2932 522356 2984
rect 524236 2932 524288 2984
rect 529020 2864 529072 2916
rect 25320 2796 25372 2848
rect 176844 2796 176896 2848
rect 182548 2796 182600 2848
rect 196716 2796 196768 2848
rect 357716 2796 357768 2848
rect 358728 2796 358780 2848
rect 359556 2796 359608 2848
rect 369400 2796 369452 2848
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 299492 703582 299980 703610
rect 8128 700330 8156 703520
rect 24320 700398 24348 703520
rect 40512 700466 40540 703520
rect 72988 700670 73016 703520
rect 89180 700738 89208 703520
rect 105464 700806 105492 703520
rect 137848 701010 137876 703520
rect 137836 701004 137888 701010
rect 137836 700946 137888 700952
rect 105452 700800 105504 700806
rect 105452 700742 105504 700748
rect 89168 700732 89220 700738
rect 89168 700674 89220 700680
rect 72976 700664 73028 700670
rect 72976 700606 73028 700612
rect 40500 700460 40552 700466
rect 40500 700402 40552 700408
rect 24308 700392 24360 700398
rect 24308 700334 24360 700340
rect 8116 700324 8168 700330
rect 8116 700266 8168 700272
rect 154132 700262 154160 703520
rect 154120 700256 154172 700262
rect 154120 700198 154172 700204
rect 170324 699718 170352 703520
rect 202800 700126 202828 703520
rect 218992 702434 219020 703520
rect 218992 702406 219388 702434
rect 202788 700120 202840 700126
rect 202788 700062 202840 700068
rect 170312 699712 170364 699718
rect 170312 699654 170364 699660
rect 171048 699712 171100 699718
rect 171048 699654 171100 699660
rect 3422 684312 3478 684321
rect 3422 684247 3478 684256
rect 3436 683194 3464 684247
rect 3424 683188 3476 683194
rect 3424 683130 3476 683136
rect 3514 671256 3570 671265
rect 3514 671191 3570 671200
rect 3528 670750 3556 671191
rect 3516 670744 3568 670750
rect 3516 670686 3568 670692
rect 3422 658200 3478 658209
rect 3422 658135 3478 658144
rect 3436 656946 3464 658135
rect 3424 656940 3476 656946
rect 3424 656882 3476 656888
rect 3424 632120 3476 632126
rect 3422 632088 3424 632097
rect 3476 632088 3478 632097
rect 3422 632023 3478 632032
rect 3146 619168 3202 619177
rect 3146 619103 3202 619112
rect 3160 618322 3188 619103
rect 3148 618316 3200 618322
rect 3148 618258 3200 618264
rect 3238 606112 3294 606121
rect 3238 606047 3294 606056
rect 3252 605878 3280 606047
rect 3240 605872 3292 605878
rect 3240 605814 3292 605820
rect 3330 580000 3386 580009
rect 3330 579935 3386 579944
rect 3344 579698 3372 579935
rect 3332 579692 3384 579698
rect 3332 579634 3384 579640
rect 3422 566944 3478 566953
rect 3422 566879 3478 566888
rect 3436 565894 3464 566879
rect 3424 565888 3476 565894
rect 3424 565830 3476 565836
rect 3422 553888 3478 553897
rect 3422 553823 3478 553832
rect 3436 553450 3464 553823
rect 3424 553444 3476 553450
rect 3424 553386 3476 553392
rect 3422 527912 3478 527921
rect 3422 527847 3478 527856
rect 3436 527202 3464 527847
rect 3424 527196 3476 527202
rect 3424 527138 3476 527144
rect 3422 514856 3478 514865
rect 3422 514791 3424 514800
rect 3476 514791 3478 514800
rect 3424 514762 3476 514768
rect 171060 511426 171088 699654
rect 219360 511494 219388 702406
rect 235184 699718 235212 703520
rect 267660 699854 267688 703520
rect 277308 700936 277360 700942
rect 277308 700878 277360 700884
rect 270408 700596 270460 700602
rect 270408 700538 270460 700544
rect 267648 699848 267700 699854
rect 267648 699790 267700 699796
rect 235172 699712 235224 699718
rect 235172 699654 235224 699660
rect 235908 699712 235960 699718
rect 235908 699654 235960 699660
rect 235920 511630 235948 699654
rect 263508 696992 263560 696998
rect 263508 696934 263560 696940
rect 260748 670812 260800 670818
rect 260748 670754 260800 670760
rect 256608 643136 256660 643142
rect 256608 643078 256660 643084
rect 255228 616888 255280 616894
rect 255228 616830 255280 616836
rect 249708 590708 249760 590714
rect 249708 590650 249760 590656
rect 248328 563100 248380 563106
rect 248328 563042 248380 563048
rect 242808 536852 242860 536858
rect 242808 536794 242860 536800
rect 235908 511624 235960 511630
rect 235908 511566 235960 511572
rect 219348 511488 219400 511494
rect 219348 511430 219400 511436
rect 171048 511420 171100 511426
rect 171048 511362 171100 511368
rect 240508 510672 240560 510678
rect 240508 510614 240560 510620
rect 198096 510604 198148 510610
rect 198096 510546 198148 510552
rect 237380 510604 237432 510610
rect 237380 510546 237432 510552
rect 238300 510604 238352 510610
rect 238300 510546 238352 510552
rect 175832 510400 175884 510406
rect 175832 510342 175884 510348
rect 100116 510196 100168 510202
rect 100116 510138 100168 510144
rect 100024 510060 100076 510066
rect 100024 510002 100076 510008
rect 82084 509924 82136 509930
rect 82084 509866 82136 509872
rect 64144 509856 64196 509862
rect 64144 509798 64196 509804
rect 4988 509720 5040 509726
rect 4988 509662 5040 509668
rect 4896 509584 4948 509590
rect 4896 509526 4948 509532
rect 4804 509312 4856 509318
rect 3422 509280 3478 509289
rect 4804 509254 4856 509260
rect 3422 509215 3478 509224
rect 3148 502308 3200 502314
rect 3148 502250 3200 502256
rect 3160 501809 3188 502250
rect 3146 501800 3202 501809
rect 3146 501735 3202 501744
rect 3332 475720 3384 475726
rect 3330 475688 3332 475697
rect 3384 475688 3386 475697
rect 3330 475623 3386 475632
rect 2780 463480 2832 463486
rect 2780 463422 2832 463428
rect 2792 462641 2820 463422
rect 2778 462632 2834 462641
rect 2778 462567 2834 462576
rect 3332 449880 3384 449886
rect 3332 449822 3384 449828
rect 3344 449585 3372 449822
rect 3330 449576 3386 449585
rect 3330 449511 3386 449520
rect 3332 423632 3384 423638
rect 3330 423600 3332 423609
rect 3384 423600 3386 423609
rect 3330 423535 3386 423544
rect 2780 411052 2832 411058
rect 2780 410994 2832 411000
rect 2792 410553 2820 410994
rect 2778 410544 2834 410553
rect 2778 410479 2834 410488
rect 3332 398812 3384 398818
rect 3332 398754 3384 398760
rect 3344 397497 3372 398754
rect 3330 397488 3386 397497
rect 3330 397423 3386 397432
rect 3056 372428 3108 372434
rect 3056 372370 3108 372376
rect 3068 371385 3096 372370
rect 3054 371376 3110 371385
rect 3054 371311 3110 371320
rect 2780 358488 2832 358494
rect 2778 358456 2780 358465
rect 2832 358456 2834 358465
rect 2778 358391 2834 358400
rect 3332 346384 3384 346390
rect 3332 346326 3384 346332
rect 3344 345409 3372 346326
rect 3330 345400 3386 345409
rect 3330 345335 3386 345344
rect 3332 319592 3384 319598
rect 3332 319534 3384 319540
rect 3344 319297 3372 319534
rect 3330 319288 3386 319297
rect 3330 319223 3386 319232
rect 3332 306332 3384 306338
rect 3332 306274 3384 306280
rect 3344 306241 3372 306274
rect 3330 306232 3386 306241
rect 3330 306167 3386 306176
rect 2872 293956 2924 293962
rect 2872 293898 2924 293904
rect 2884 293185 2912 293898
rect 2870 293176 2926 293185
rect 2870 293111 2926 293120
rect 3240 267708 3292 267714
rect 3240 267650 3292 267656
rect 3252 267209 3280 267650
rect 3238 267200 3294 267209
rect 3238 267135 3294 267144
rect 3332 255264 3384 255270
rect 3332 255206 3384 255212
rect 3344 254153 3372 255206
rect 3330 254144 3386 254153
rect 3330 254079 3386 254088
rect 3332 215008 3384 215014
rect 3330 214976 3332 214985
rect 3384 214976 3386 214985
rect 3330 214911 3386 214920
rect 3056 202836 3108 202842
rect 3056 202778 3108 202784
rect 3068 201929 3096 202778
rect 3054 201920 3110 201929
rect 3054 201855 3110 201864
rect 2780 188896 2832 188902
rect 2778 188864 2780 188873
rect 2832 188864 2834 188873
rect 2778 188799 2834 188808
rect 3332 164212 3384 164218
rect 3332 164154 3384 164160
rect 3344 162897 3372 164154
rect 3330 162888 3386 162897
rect 3330 162823 3386 162832
rect 3056 59356 3108 59362
rect 3056 59298 3108 59304
rect 3068 58585 3096 59298
rect 3054 58576 3110 58585
rect 3054 58511 3110 58520
rect 2872 33108 2924 33114
rect 2872 33050 2924 33056
rect 2884 32473 2912 33050
rect 2870 32464 2926 32473
rect 2870 32399 2926 32408
rect 3436 6497 3464 509215
rect 3608 506592 3660 506598
rect 3608 506534 3660 506540
rect 3516 506524 3568 506530
rect 3516 506466 3568 506472
rect 3528 136785 3556 506466
rect 3620 241097 3648 506534
rect 3606 241088 3662 241097
rect 3606 241023 3662 241032
rect 4816 188902 4844 509254
rect 4908 358494 4936 509526
rect 5000 411058 5028 509662
rect 14648 509652 14700 509658
rect 14648 509594 14700 509600
rect 11704 509516 11756 509522
rect 11704 509458 11756 509464
rect 7932 508564 7984 508570
rect 7932 508506 7984 508512
rect 7840 508496 7892 508502
rect 7840 508438 7892 508444
rect 7748 508360 7800 508366
rect 7748 508302 7800 508308
rect 7656 508020 7708 508026
rect 7656 507962 7708 507968
rect 7564 507952 7616 507958
rect 7564 507894 7616 507900
rect 5540 507068 5592 507074
rect 5540 507010 5592 507016
rect 5080 506864 5132 506870
rect 5080 506806 5132 506812
rect 5092 463486 5120 506806
rect 5552 502314 5580 507010
rect 5540 502308 5592 502314
rect 5540 502250 5592 502256
rect 5080 463480 5132 463486
rect 5080 463422 5132 463428
rect 4988 411052 5040 411058
rect 4988 410994 5040 411000
rect 4896 358488 4948 358494
rect 4896 358430 4948 358436
rect 4804 188896 4856 188902
rect 4804 188838 4856 188844
rect 3608 150408 3660 150414
rect 3608 150350 3660 150356
rect 3620 149841 3648 150350
rect 3606 149832 3662 149841
rect 3606 149767 3662 149776
rect 3514 136776 3570 136785
rect 3514 136711 3570 136720
rect 3516 110764 3568 110770
rect 3516 110706 3568 110712
rect 3528 110673 3556 110706
rect 3514 110664 3570 110673
rect 3514 110599 3570 110608
rect 3516 97980 3568 97986
rect 3516 97922 3568 97928
rect 3528 97617 3556 97922
rect 3514 97608 3570 97617
rect 3514 97543 3570 97552
rect 3516 85536 3568 85542
rect 3516 85478 3568 85484
rect 3528 84697 3556 85478
rect 3514 84688 3570 84697
rect 3514 84623 3570 84632
rect 7576 71670 7604 507894
rect 7668 110770 7696 507962
rect 7760 372434 7788 508302
rect 7852 423638 7880 508438
rect 7944 475726 7972 508506
rect 9036 508292 9088 508298
rect 9036 508234 9088 508240
rect 8944 508156 8996 508162
rect 8944 508098 8996 508104
rect 7932 475720 7984 475726
rect 7932 475662 7984 475668
rect 7840 423632 7892 423638
rect 7840 423574 7892 423580
rect 7748 372428 7800 372434
rect 7748 372370 7800 372376
rect 8956 215014 8984 508098
rect 9048 319598 9076 508234
rect 10508 508224 10560 508230
rect 10508 508166 10560 508172
rect 10416 508088 10468 508094
rect 10416 508030 10468 508036
rect 10324 507884 10376 507890
rect 10324 507826 10376 507832
rect 9036 319592 9088 319598
rect 9036 319534 9088 319540
rect 8944 215008 8996 215014
rect 8944 214950 8996 214956
rect 7656 110764 7708 110770
rect 7656 110706 7708 110712
rect 3516 71664 3568 71670
rect 3514 71632 3516 71641
rect 7564 71664 7616 71670
rect 3568 71632 3570 71641
rect 7564 71606 7616 71612
rect 3514 71567 3570 71576
rect 3516 45552 3568 45558
rect 3514 45520 3516 45529
rect 3568 45520 3570 45529
rect 3514 45455 3570 45464
rect 10336 33114 10364 507826
rect 10428 164218 10456 508030
rect 10520 267714 10548 508166
rect 11716 306338 11744 509458
rect 14556 509448 14608 509454
rect 14556 509390 14608 509396
rect 14464 509380 14516 509386
rect 14464 509322 14516 509328
rect 11980 507000 12032 507006
rect 11980 506942 12032 506948
rect 11888 506932 11940 506938
rect 11888 506874 11940 506880
rect 11796 506796 11848 506802
rect 11796 506738 11848 506744
rect 11808 346390 11836 506738
rect 11900 398818 11928 506874
rect 11992 449886 12020 506942
rect 11980 449880 12032 449886
rect 11980 449822 12032 449828
rect 11888 398812 11940 398818
rect 11888 398754 11940 398760
rect 11796 346384 11848 346390
rect 11796 346326 11848 346332
rect 11704 306332 11756 306338
rect 11704 306274 11756 306280
rect 10508 267708 10560 267714
rect 10508 267650 10560 267656
rect 14476 202842 14504 509322
rect 14568 255270 14596 509390
rect 14660 293962 14688 509594
rect 14648 293956 14700 293962
rect 14648 293898 14700 293904
rect 14556 255264 14608 255270
rect 14556 255206 14608 255212
rect 14464 202836 14516 202842
rect 14464 202778 14516 202784
rect 61384 198688 61436 198694
rect 61384 198630 61436 198636
rect 58624 198484 58676 198490
rect 58624 198426 58676 198432
rect 51724 198416 51776 198422
rect 51724 198358 51776 198364
rect 35164 198280 35216 198286
rect 35164 198222 35216 198228
rect 29644 198212 29696 198218
rect 29644 198154 29696 198160
rect 18604 198144 18656 198150
rect 18604 198086 18656 198092
rect 11704 198076 11756 198082
rect 11704 198018 11756 198024
rect 10416 164212 10468 164218
rect 10416 164154 10468 164160
rect 10324 33108 10376 33114
rect 10324 33050 10376 33056
rect 3516 20664 3568 20670
rect 3516 20606 3568 20612
rect 3528 19417 3556 20606
rect 3514 19408 3570 19417
rect 3514 19343 3570 19352
rect 3422 6488 3478 6497
rect 3422 6423 3478 6432
rect 8760 6248 8812 6254
rect 8760 6190 8812 6196
rect 4068 6180 4120 6186
rect 4068 6122 4120 6128
rect 2872 4956 2924 4962
rect 2872 4898 2924 4904
rect 1676 4888 1728 4894
rect 1676 4830 1728 4836
rect 572 4820 624 4826
rect 572 4762 624 4768
rect 584 480 612 4762
rect 1688 480 1716 4830
rect 2884 480 2912 4898
rect 4080 480 4108 6122
rect 7656 5024 7708 5030
rect 7656 4966 7708 4972
rect 5264 3528 5316 3534
rect 5264 3470 5316 3476
rect 5276 480 5304 3470
rect 6460 3460 6512 3466
rect 6460 3402 6512 3408
rect 6472 480 6500 3402
rect 7668 480 7696 4966
rect 8772 480 8800 6190
rect 11152 4072 11204 4078
rect 11152 4014 11204 4020
rect 9956 3256 10008 3262
rect 9956 3198 10008 3204
rect 9968 480 9996 3198
rect 11164 480 11192 4014
rect 11716 3534 11744 198018
rect 14464 198008 14516 198014
rect 14464 197950 14516 197956
rect 12348 5092 12400 5098
rect 12348 5034 12400 5040
rect 11704 3528 11756 3534
rect 11704 3470 11756 3476
rect 12360 480 12388 5034
rect 13544 3528 13596 3534
rect 13544 3470 13596 3476
rect 13556 480 13584 3470
rect 14476 3262 14504 197950
rect 14556 196648 14608 196654
rect 14556 196590 14608 196596
rect 14568 3534 14596 196590
rect 17040 4208 17092 4214
rect 17040 4150 17092 4156
rect 15936 3596 15988 3602
rect 15936 3538 15988 3544
rect 14556 3528 14608 3534
rect 14556 3470 14608 3476
rect 14740 3528 14792 3534
rect 14740 3470 14792 3476
rect 14464 3256 14516 3262
rect 14464 3198 14516 3204
rect 14752 480 14780 3470
rect 15948 480 15976 3538
rect 17052 480 17080 4150
rect 18616 4078 18644 198086
rect 23388 89004 23440 89010
rect 23388 88946 23440 88952
rect 19248 14476 19300 14482
rect 19248 14418 19300 14424
rect 18604 4072 18656 4078
rect 18604 4014 18656 4020
rect 19260 3398 19288 14418
rect 23400 6914 23428 88946
rect 28908 87644 28960 87650
rect 28908 87586 28960 87592
rect 23032 6886 23428 6914
rect 21824 6316 21876 6322
rect 21824 6258 21876 6264
rect 20628 4072 20680 4078
rect 20628 4014 20680 4020
rect 19432 3800 19484 3806
rect 19432 3742 19484 3748
rect 18236 3392 18288 3398
rect 18236 3334 18288 3340
rect 19248 3392 19300 3398
rect 19248 3334 19300 3340
rect 18248 480 18276 3334
rect 19444 480 19472 3742
rect 20640 480 20668 4014
rect 21836 480 21864 6258
rect 23032 480 23060 6886
rect 26516 6384 26568 6390
rect 26516 6326 26568 6332
rect 24216 3664 24268 3670
rect 24216 3606 24268 3612
rect 24228 480 24256 3606
rect 25320 2848 25372 2854
rect 25320 2790 25372 2796
rect 25332 480 25360 2790
rect 26528 480 26556 6326
rect 28920 3398 28948 87586
rect 29656 3806 29684 198154
rect 32404 22772 32456 22778
rect 32404 22714 32456 22720
rect 30104 6452 30156 6458
rect 30104 6394 30156 6400
rect 29644 3800 29696 3806
rect 29644 3742 29696 3748
rect 27712 3392 27764 3398
rect 27712 3334 27764 3340
rect 28908 3392 28960 3398
rect 28908 3334 28960 3340
rect 27724 480 27752 3334
rect 28908 3256 28960 3262
rect 28908 3198 28960 3204
rect 28920 480 28948 3198
rect 30116 480 30144 6394
rect 32416 3398 32444 22714
rect 33600 6520 33652 6526
rect 33600 6462 33652 6468
rect 32496 3800 32548 3806
rect 32496 3742 32548 3748
rect 31300 3392 31352 3398
rect 31300 3334 31352 3340
rect 32404 3392 32456 3398
rect 32404 3334 32456 3340
rect 31312 480 31340 3334
rect 32508 1986 32536 3742
rect 32416 1958 32536 1986
rect 32416 480 32444 1958
rect 33612 480 33640 6462
rect 34796 3392 34848 3398
rect 34796 3334 34848 3340
rect 34808 480 34836 3334
rect 35176 3262 35204 198222
rect 39304 196716 39356 196722
rect 39304 196658 39356 196664
rect 35808 89072 35860 89078
rect 35808 89014 35860 89020
rect 35820 3398 35848 89014
rect 37188 6588 37240 6594
rect 37188 6530 37240 6536
rect 35992 4072 36044 4078
rect 35992 4014 36044 4020
rect 35808 3392 35860 3398
rect 35808 3334 35860 3340
rect 35164 3256 35216 3262
rect 35164 3198 35216 3204
rect 36004 480 36032 4014
rect 37200 480 37228 6530
rect 39316 3398 39344 196658
rect 43444 87712 43496 87718
rect 43444 87654 43496 87660
rect 40684 6656 40736 6662
rect 40684 6598 40736 6604
rect 39580 3868 39632 3874
rect 39580 3810 39632 3816
rect 38384 3392 38436 3398
rect 38384 3334 38436 3340
rect 39304 3392 39356 3398
rect 39304 3334 39356 3340
rect 38396 480 38424 3334
rect 39592 480 39620 3810
rect 40696 480 40724 6598
rect 43456 3398 43484 87654
rect 45468 15904 45520 15910
rect 45468 15846 45520 15852
rect 44272 6724 44324 6730
rect 44272 6666 44324 6672
rect 41880 3392 41932 3398
rect 41880 3334 41932 3340
rect 43444 3392 43496 3398
rect 43444 3334 43496 3340
rect 41892 480 41920 3334
rect 43076 3324 43128 3330
rect 43076 3266 43128 3272
rect 43088 480 43116 3266
rect 44284 480 44312 6666
rect 45480 480 45508 15846
rect 48964 7608 49016 7614
rect 48964 7550 49016 7556
rect 47860 5228 47912 5234
rect 47860 5170 47912 5176
rect 46664 3936 46716 3942
rect 46664 3878 46716 3884
rect 46676 480 46704 3878
rect 47872 480 47900 5170
rect 48976 480 49004 7550
rect 51356 5296 51408 5302
rect 51356 5238 51408 5244
rect 50160 4004 50212 4010
rect 50160 3946 50212 3952
rect 50172 480 50200 3946
rect 51368 480 51396 5238
rect 51736 4078 51764 198358
rect 57244 198348 57296 198354
rect 57244 198290 57296 198296
rect 56048 7744 56100 7750
rect 56048 7686 56100 7692
rect 52552 7676 52604 7682
rect 52552 7618 52604 7624
rect 51724 4072 51776 4078
rect 51724 4014 51776 4020
rect 52564 480 52592 7618
rect 54944 5364 54996 5370
rect 54944 5306 54996 5312
rect 53748 4072 53800 4078
rect 53748 4014 53800 4020
rect 53760 480 53788 4014
rect 54956 480 54984 5306
rect 56060 480 56088 7686
rect 57256 6914 57284 198290
rect 57164 6886 57284 6914
rect 57164 4078 57192 6886
rect 58440 5432 58492 5438
rect 58440 5374 58492 5380
rect 57152 4072 57204 4078
rect 57152 4014 57204 4020
rect 57244 4072 57296 4078
rect 57244 4014 57296 4020
rect 57256 480 57284 4014
rect 58452 480 58480 5374
rect 58636 3398 58664 198426
rect 59636 7812 59688 7818
rect 59636 7754 59688 7760
rect 58624 3392 58676 3398
rect 58624 3334 58676 3340
rect 59648 480 59676 7754
rect 61396 4146 61424 198630
rect 64156 85542 64184 509798
rect 76564 198620 76616 198626
rect 76564 198562 76616 198568
rect 71044 198552 71096 198558
rect 71044 198494 71096 198500
rect 64144 85536 64196 85542
rect 64144 85478 64196 85484
rect 70308 9104 70360 9110
rect 70308 9046 70360 9052
rect 66720 9036 66772 9042
rect 66720 8978 66772 8984
rect 63224 8968 63276 8974
rect 63224 8910 63276 8916
rect 62028 5500 62080 5506
rect 62028 5442 62080 5448
rect 61384 4140 61436 4146
rect 61384 4082 61436 4088
rect 60832 3324 60884 3330
rect 60832 3266 60884 3272
rect 60844 480 60872 3266
rect 62040 480 62068 5442
rect 63236 480 63264 8910
rect 65524 4752 65576 4758
rect 65524 4694 65576 4700
rect 64328 4140 64380 4146
rect 64328 4082 64380 4088
rect 64340 480 64368 4082
rect 65536 480 65564 4694
rect 66732 480 66760 8978
rect 69112 4616 69164 4622
rect 69112 4558 69164 4564
rect 67916 3732 67968 3738
rect 67916 3674 67968 3680
rect 67928 480 67956 3674
rect 69124 480 69152 4558
rect 70320 480 70348 9046
rect 71056 3330 71084 198494
rect 73804 9172 73856 9178
rect 73804 9114 73856 9120
rect 72608 4684 72660 4690
rect 72608 4626 72660 4632
rect 71504 3392 71556 3398
rect 71504 3334 71556 3340
rect 71044 3324 71096 3330
rect 71044 3266 71096 3272
rect 71516 480 71544 3334
rect 72620 480 72648 4626
rect 73816 480 73844 9114
rect 76196 4548 76248 4554
rect 76196 4490 76248 4496
rect 75000 3120 75052 3126
rect 75000 3062 75052 3068
rect 75012 480 75040 3062
rect 76208 480 76236 4490
rect 76576 3738 76604 198562
rect 81348 89140 81400 89146
rect 81348 89082 81400 89088
rect 77392 9240 77444 9246
rect 77392 9182 77444 9188
rect 76564 3732 76616 3738
rect 76564 3674 76616 3680
rect 77404 480 77432 9182
rect 79692 6792 79744 6798
rect 79692 6734 79744 6740
rect 78588 3324 78640 3330
rect 78588 3266 78640 3272
rect 78600 480 78628 3266
rect 79704 480 79732 6734
rect 81360 3738 81388 89082
rect 82096 45558 82124 509866
rect 94504 197940 94556 197946
rect 94504 197882 94556 197888
rect 88248 196784 88300 196790
rect 88248 196726 88300 196732
rect 82084 45552 82136 45558
rect 82084 45494 82136 45500
rect 85488 14544 85540 14550
rect 85488 14486 85540 14492
rect 83280 6860 83332 6866
rect 83280 6802 83332 6808
rect 80888 3732 80940 3738
rect 80888 3674 80940 3680
rect 81348 3732 81400 3738
rect 81348 3674 81400 3680
rect 80900 480 80928 3674
rect 82084 3052 82136 3058
rect 82084 2994 82136 3000
rect 82096 480 82124 2994
rect 83292 480 83320 6802
rect 85500 3738 85528 14486
rect 86868 7880 86920 7886
rect 86868 7822 86920 7828
rect 84476 3732 84528 3738
rect 84476 3674 84528 3680
rect 85488 3732 85540 3738
rect 85488 3674 85540 3680
rect 84488 480 84516 3674
rect 85672 2984 85724 2990
rect 85672 2926 85724 2932
rect 85684 480 85712 2926
rect 86880 480 86908 7822
rect 88260 6914 88288 196726
rect 92388 15972 92440 15978
rect 92388 15914 92440 15920
rect 90364 7948 90416 7954
rect 90364 7890 90416 7896
rect 87984 6886 88288 6914
rect 87984 480 88012 6886
rect 89168 3256 89220 3262
rect 89168 3198 89220 3204
rect 89180 480 89208 3198
rect 90376 480 90404 7890
rect 92400 3738 92428 15914
rect 93952 8016 94004 8022
rect 93952 7958 94004 7964
rect 91560 3732 91612 3738
rect 91560 3674 91612 3680
rect 92388 3732 92440 3738
rect 92388 3674 92440 3680
rect 92756 3732 92808 3738
rect 92756 3674 92808 3680
rect 91572 480 91600 3674
rect 92768 480 92796 3674
rect 93964 480 93992 7958
rect 94516 3738 94544 197882
rect 98644 197668 98696 197674
rect 98644 197610 98696 197616
rect 95148 84856 95200 84862
rect 95148 84798 95200 84804
rect 94504 3732 94556 3738
rect 94504 3674 94556 3680
rect 95160 480 95188 84798
rect 97448 8084 97500 8090
rect 97448 8026 97500 8032
rect 96252 3188 96304 3194
rect 96252 3130 96304 3136
rect 96264 480 96292 3130
rect 97460 480 97488 8026
rect 98656 6914 98684 197610
rect 100036 59362 100064 510002
rect 100128 150414 100156 510138
rect 101496 510128 101548 510134
rect 101496 510070 101548 510076
rect 101404 509992 101456 509998
rect 101404 509934 101456 509940
rect 100116 150408 100168 150414
rect 100116 150350 100168 150356
rect 100024 59356 100076 59362
rect 100024 59298 100076 59304
rect 99288 44872 99340 44878
rect 99288 44814 99340 44820
rect 98564 6886 98684 6914
rect 98564 3126 98592 6886
rect 99300 3738 99328 44814
rect 101416 20670 101444 509934
rect 101508 97986 101536 510070
rect 173532 508700 173584 508706
rect 173532 508642 173584 508648
rect 169116 508632 169168 508638
rect 169116 508574 169168 508580
rect 166814 507920 166870 507929
rect 166870 507878 166934 507906
rect 169128 507892 169156 508574
rect 173544 507892 173572 508642
rect 175844 507892 175872 510342
rect 193680 508904 193732 508910
rect 193680 508846 193732 508852
rect 186964 508836 187016 508842
rect 186964 508778 187016 508784
rect 180248 508768 180300 508774
rect 180248 508710 180300 508716
rect 180260 507892 180288 508710
rect 186976 507892 187004 508778
rect 193692 507892 193720 508846
rect 198108 507892 198136 510546
rect 231584 510536 231636 510542
rect 231584 510478 231636 510484
rect 229376 510468 229428 510474
rect 229376 510410 229428 510416
rect 215944 510332 215996 510338
rect 215944 510274 215996 510280
rect 213736 509108 213788 509114
rect 213736 509050 213788 509056
rect 207020 509040 207072 509046
rect 207020 508982 207072 508988
rect 200396 508972 200448 508978
rect 200396 508914 200448 508920
rect 200408 507892 200436 508914
rect 207032 507892 207060 508982
rect 213748 507892 213776 509050
rect 215956 507892 215984 510274
rect 224960 510264 225012 510270
rect 224960 510206 225012 510212
rect 222660 509788 222712 509794
rect 222660 509730 222712 509736
rect 220452 508428 220504 508434
rect 220452 508370 220504 508376
rect 220464 507892 220492 508370
rect 222672 507892 222700 509730
rect 224972 507892 225000 510206
rect 229388 507892 229416 510410
rect 231596 507892 231624 510478
rect 237392 509250 237420 510546
rect 237380 509244 237432 509250
rect 237380 509186 237432 509192
rect 233884 509176 233936 509182
rect 233884 509118 233936 509124
rect 233896 507892 233924 509118
rect 238312 507892 238340 510546
rect 240520 507892 240548 510614
rect 242820 507892 242848 536794
rect 245568 524476 245620 524482
rect 245568 524418 245620 524424
rect 245580 509234 245608 524418
rect 248340 509234 248368 563042
rect 245488 509206 245608 509234
rect 247696 509206 248368 509234
rect 245488 507906 245516 509206
rect 247696 507906 247724 509206
rect 249720 507906 249748 590650
rect 252468 576904 252520 576910
rect 252468 576846 252520 576852
rect 252480 509234 252508 576846
rect 255240 509234 255268 616830
rect 256620 509234 256648 643078
rect 259368 630692 259420 630698
rect 259368 630634 259420 630640
rect 259380 509234 259408 630634
rect 252112 509206 252508 509234
rect 254320 509206 255268 509234
rect 256528 509206 256648 509234
rect 258920 509206 259408 509234
rect 252112 507906 252140 509206
rect 254320 507906 254348 509206
rect 256528 507906 256556 509206
rect 258920 507906 258948 509206
rect 260760 507906 260788 670754
rect 263520 509234 263548 696934
rect 266268 683256 266320 683262
rect 266268 683198 266320 683204
rect 266280 509234 266308 683198
rect 267372 511284 267424 511290
rect 267372 511226 267424 511232
rect 263336 509206 263548 509234
rect 265544 509206 266308 509234
rect 263336 507906 263364 509206
rect 265544 507906 265572 509206
rect 245042 507878 245516 507906
rect 247250 507878 247724 507906
rect 249550 507878 249748 507906
rect 251758 507878 252140 507906
rect 253966 507878 254348 507906
rect 256174 507878 256556 507906
rect 258474 507878 258948 507906
rect 260682 507878 260788 507906
rect 262890 507878 263364 507906
rect 265098 507878 265572 507906
rect 267384 507892 267412 511226
rect 270420 509234 270448 700538
rect 271788 700528 271840 700534
rect 271788 700470 271840 700476
rect 269960 509206 270448 509234
rect 269960 507906 269988 509206
rect 269606 507878 269988 507906
rect 271800 507892 271828 700470
rect 274088 511352 274140 511358
rect 274088 511294 274140 511300
rect 274100 507892 274128 511294
rect 277320 509234 277348 700878
rect 278688 700868 278740 700874
rect 278688 700810 278740 700816
rect 276768 509206 277348 509234
rect 276768 507906 276796 509206
rect 278700 507906 278728 700810
rect 283852 699786 283880 703520
rect 285588 700188 285640 700194
rect 285588 700130 285640 700136
rect 284208 700052 284260 700058
rect 284208 699994 284260 700000
rect 283840 699780 283892 699786
rect 283840 699722 283892 699728
rect 280712 511692 280764 511698
rect 280712 511634 280764 511640
rect 276322 507878 276796 507906
rect 278530 507878 278728 507906
rect 280724 507892 280752 511634
rect 284220 509234 284248 699994
rect 283392 509206 284248 509234
rect 283392 507906 283420 509206
rect 285600 507906 285628 700130
rect 292488 699984 292540 699990
rect 292488 699926 292540 699932
rect 289728 699916 289780 699922
rect 289728 699858 289780 699864
rect 287428 511556 287480 511562
rect 287428 511498 287480 511504
rect 283038 507878 283420 507906
rect 285246 507878 285628 507906
rect 287440 507892 287468 511498
rect 289740 507906 289768 699858
rect 292500 509234 292528 699926
rect 295340 699848 295392 699854
rect 295340 699790 295392 699796
rect 295352 518894 295380 699790
rect 298100 699780 298152 699786
rect 298100 699722 298152 699728
rect 298112 518894 298140 699722
rect 295352 518866 296024 518894
rect 298112 518866 298232 518894
rect 294144 511760 294196 511766
rect 294144 511702 294196 511708
rect 292408 509206 292528 509234
rect 292408 507906 292436 509206
rect 289662 507878 289768 507906
rect 291962 507878 292436 507906
rect 294156 507892 294184 511702
rect 295996 507906 296024 518866
rect 298204 507906 298232 518866
rect 299492 511766 299520 703582
rect 299952 703474 299980 703582
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494072 703582 494652 703610
rect 300136 703474 300164 703520
rect 299952 703446 300164 703474
rect 309140 701004 309192 701010
rect 309140 700946 309192 700952
rect 302240 700120 302292 700126
rect 302240 700062 302292 700068
rect 302884 700120 302936 700126
rect 302884 700062 302936 700068
rect 302252 518894 302280 700062
rect 302252 518866 302648 518894
rect 299480 511760 299532 511766
rect 299480 511702 299532 511708
rect 300860 511624 300912 511630
rect 300860 511566 300912 511572
rect 295996 507878 296378 507906
rect 298204 507878 298678 507906
rect 300872 507892 300900 511566
rect 302620 507906 302648 518866
rect 302896 511698 302924 700062
rect 309152 518894 309180 700946
rect 313280 700800 313332 700806
rect 313280 700742 313332 700748
rect 311900 700256 311952 700262
rect 311900 700198 311952 700204
rect 309152 518866 309456 518894
rect 302884 511692 302936 511698
rect 302884 511634 302936 511640
rect 305276 511488 305328 511494
rect 305276 511430 305328 511436
rect 302620 507878 303094 507906
rect 305288 507892 305316 511430
rect 307576 511420 307628 511426
rect 307576 511362 307628 511368
rect 307588 507892 307616 511362
rect 309428 507906 309456 518866
rect 311912 507906 311940 700198
rect 313292 518894 313320 700742
rect 317420 700732 317472 700738
rect 317420 700674 317472 700680
rect 316040 700664 316092 700670
rect 316040 700606 316092 700612
rect 313292 518866 313872 518894
rect 313844 507906 313872 518866
rect 316052 507906 316080 700606
rect 317432 518894 317460 700674
rect 320180 700460 320232 700466
rect 320180 700402 320232 700408
rect 320192 518894 320220 700402
rect 324320 700392 324372 700398
rect 324320 700334 324372 700340
rect 322940 700324 322992 700330
rect 322940 700266 322992 700272
rect 317432 518866 318288 518894
rect 320192 518866 320496 518894
rect 318260 507906 318288 518866
rect 320468 507906 320496 518866
rect 322952 507906 322980 700266
rect 324332 518894 324360 700334
rect 332520 699922 332548 703520
rect 348804 699990 348832 703520
rect 364996 702434 365024 703520
rect 364352 702406 365024 702434
rect 348792 699984 348844 699990
rect 348792 699926 348844 699932
rect 332508 699916 332560 699922
rect 332508 699858 332560 699864
rect 327080 683188 327132 683194
rect 327080 683130 327132 683136
rect 327092 518894 327120 683130
rect 331220 670744 331272 670750
rect 331220 670686 331272 670692
rect 329840 656940 329892 656946
rect 329840 656882 329892 656888
rect 324332 518866 325096 518894
rect 327092 518866 327304 518894
rect 325068 507906 325096 518866
rect 327276 507906 327304 518866
rect 309428 507878 309810 507906
rect 311912 507878 312018 507906
rect 313844 507878 314226 507906
rect 316052 507878 316526 507906
rect 318260 507878 318734 507906
rect 320468 507878 320942 507906
rect 322952 507878 323242 507906
rect 325068 507878 325450 507906
rect 327276 507878 327658 507906
rect 329852 507892 329880 656882
rect 331232 518894 331260 670686
rect 333980 632120 334032 632126
rect 333980 632062 334032 632068
rect 331232 518866 331720 518894
rect 331692 507906 331720 518866
rect 333992 507906 334020 632062
rect 338120 618316 338172 618322
rect 338120 618258 338172 618264
rect 335360 605872 335412 605878
rect 335360 605814 335412 605820
rect 335372 518894 335400 605814
rect 338132 518894 338160 618258
rect 340880 579692 340932 579698
rect 340880 579634 340932 579640
rect 335372 518866 336136 518894
rect 338132 518866 338344 518894
rect 336108 507906 336136 518866
rect 338316 507906 338344 518866
rect 340892 507906 340920 579634
rect 345020 565888 345072 565894
rect 345020 565830 345072 565836
rect 342260 553444 342312 553450
rect 342260 553386 342312 553392
rect 342272 518894 342300 553386
rect 345032 518894 345060 565830
rect 347780 527196 347832 527202
rect 347780 527138 347832 527144
rect 342272 518866 342944 518894
rect 345032 518866 345152 518894
rect 342916 507906 342944 518866
rect 345124 507906 345152 518866
rect 331692 507878 332166 507906
rect 333992 507878 334374 507906
rect 336108 507878 336582 507906
rect 338316 507878 338790 507906
rect 340892 507878 341090 507906
rect 342916 507878 343298 507906
rect 345124 507878 345506 507906
rect 347792 507892 347820 527138
rect 351920 514820 351972 514826
rect 351920 514762 351972 514768
rect 351932 507906 351960 514762
rect 364352 511562 364380 702406
rect 397472 700058 397500 703520
rect 413664 700194 413692 703520
rect 413652 700188 413704 700194
rect 413652 700130 413704 700136
rect 429856 700126 429884 703520
rect 462332 700942 462360 703520
rect 462320 700936 462372 700942
rect 462320 700878 462372 700884
rect 478524 700874 478552 703520
rect 478512 700868 478564 700874
rect 478512 700810 478564 700816
rect 429844 700120 429896 700126
rect 429844 700062 429896 700068
rect 397460 700052 397512 700058
rect 397460 699994 397512 700000
rect 364340 511556 364392 511562
rect 364340 511498 364392 511504
rect 494072 511358 494100 703582
rect 494624 703474 494652 703582
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 494808 703474 494836 703520
rect 494624 703446 494836 703474
rect 527192 700602 527220 703520
rect 527180 700596 527232 700602
rect 527180 700538 527232 700544
rect 543476 700534 543504 703520
rect 559668 702434 559696 703520
rect 558932 702406 559696 702434
rect 543464 700528 543516 700534
rect 543464 700470 543516 700476
rect 494060 511352 494112 511358
rect 494060 511294 494112 511300
rect 558932 511290 558960 702406
rect 580170 697232 580226 697241
rect 580170 697167 580226 697176
rect 580184 696998 580212 697167
rect 580172 696992 580224 696998
rect 580172 696934 580224 696940
rect 580170 683904 580226 683913
rect 580170 683839 580226 683848
rect 580184 683262 580212 683839
rect 580172 683256 580224 683262
rect 580172 683198 580224 683204
rect 580172 670812 580224 670818
rect 580172 670754 580224 670760
rect 580184 670721 580212 670754
rect 580170 670712 580226 670721
rect 580170 670647 580226 670656
rect 580170 644056 580226 644065
rect 580170 643991 580226 644000
rect 580184 643142 580212 643991
rect 580172 643136 580224 643142
rect 580172 643078 580224 643084
rect 580170 630864 580226 630873
rect 580170 630799 580226 630808
rect 580184 630698 580212 630799
rect 580172 630692 580224 630698
rect 580172 630634 580224 630640
rect 580170 617536 580226 617545
rect 580170 617471 580226 617480
rect 580184 616894 580212 617471
rect 580172 616888 580224 616894
rect 580172 616830 580224 616836
rect 579802 591016 579858 591025
rect 579802 590951 579858 590960
rect 579816 590714 579844 590951
rect 579804 590708 579856 590714
rect 579804 590650 579856 590656
rect 580170 577688 580226 577697
rect 580170 577623 580226 577632
rect 580184 576910 580212 577623
rect 580172 576904 580224 576910
rect 580172 576846 580224 576852
rect 579802 564360 579858 564369
rect 579802 564295 579858 564304
rect 579816 563106 579844 564295
rect 579804 563100 579856 563106
rect 579804 563042 579856 563048
rect 580170 537840 580226 537849
rect 580170 537775 580226 537784
rect 580184 536858 580212 537775
rect 580172 536852 580224 536858
rect 580172 536794 580224 536800
rect 580170 524512 580226 524521
rect 580170 524447 580172 524456
rect 580224 524447 580226 524456
rect 580172 524418 580224 524424
rect 580170 511320 580226 511329
rect 558920 511284 558972 511290
rect 580170 511255 580226 511264
rect 558920 511226 558972 511232
rect 580184 510678 580212 511255
rect 580172 510672 580224 510678
rect 580172 510614 580224 510620
rect 431316 510604 431368 510610
rect 431316 510546 431368 510552
rect 431224 510536 431276 510542
rect 431224 510478 431276 510484
rect 430120 510468 430172 510474
rect 430120 510410 430172 510416
rect 424324 510400 424376 510406
rect 424324 510342 424376 510348
rect 399116 510196 399168 510202
rect 399116 510138 399168 510144
rect 365628 509720 365680 509726
rect 365628 509662 365680 509668
rect 354404 508564 354456 508570
rect 354404 508506 354456 508512
rect 361120 508564 361172 508570
rect 361120 508506 361172 508512
rect 351932 507878 352222 507906
rect 354416 507892 354444 508506
rect 356704 508496 356756 508502
rect 356704 508438 356756 508444
rect 358912 508496 358964 508502
rect 358912 508438 358964 508444
rect 356716 507892 356744 508438
rect 358924 507892 358952 508438
rect 361132 507892 361160 508506
rect 363328 508496 363380 508502
rect 363328 508438 363380 508444
rect 363340 507892 363368 508438
rect 365640 507892 365668 509662
rect 376760 509652 376812 509658
rect 376760 509594 376812 509600
rect 372344 509584 372396 509590
rect 372344 509526 372396 509532
rect 367836 508360 367888 508366
rect 367836 508302 367888 508308
rect 370044 508360 370096 508366
rect 370044 508302 370096 508308
rect 367848 507892 367876 508302
rect 370056 507892 370084 508302
rect 372356 507892 372384 509526
rect 374552 508292 374604 508298
rect 374552 508234 374604 508240
rect 374564 507892 374592 508234
rect 376772 507892 376800 509594
rect 378968 509516 379020 509522
rect 378968 509458 379020 509464
rect 378980 507892 379008 509458
rect 385684 509448 385736 509454
rect 385684 509390 385736 509396
rect 381268 508224 381320 508230
rect 381268 508166 381320 508172
rect 383476 508224 383528 508230
rect 383476 508166 383528 508172
rect 381280 507892 381308 508166
rect 383488 507892 383516 508166
rect 385696 507892 385724 509390
rect 392400 509380 392452 509386
rect 392400 509322 392452 509328
rect 390192 509312 390244 509318
rect 390192 509254 390244 509260
rect 387892 508156 387944 508162
rect 387892 508098 387944 508104
rect 387904 507892 387932 508098
rect 390204 507892 390232 509254
rect 392412 507892 392440 509322
rect 394608 508088 394660 508094
rect 394608 508030 394660 508036
rect 394620 507892 394648 508030
rect 396540 508020 396592 508026
rect 396540 507962 396592 507968
rect 396552 507906 396580 507962
rect 396552 507878 396934 507906
rect 399128 507892 399156 510138
rect 405832 510128 405884 510134
rect 405832 510070 405884 510076
rect 403532 509856 403584 509862
rect 403532 509798 403584 509804
rect 401324 508088 401376 508094
rect 401324 508030 401376 508036
rect 401336 507892 401364 508030
rect 403544 507892 403572 509798
rect 405844 507892 405872 510070
rect 412456 510060 412508 510066
rect 412456 510002 412508 510008
rect 410248 509924 410300 509930
rect 410248 509866 410300 509872
rect 407764 507952 407816 507958
rect 407816 507900 408066 507906
rect 407764 507894 408066 507900
rect 407776 507878 408066 507894
rect 410260 507892 410288 509866
rect 412468 507892 412496 510002
rect 419172 509992 419224 509998
rect 419172 509934 419224 509940
rect 416962 509280 417018 509289
rect 416962 509215 417018 509224
rect 414400 507890 414782 507906
rect 416976 507892 417004 509215
rect 419184 507892 419212 509934
rect 421932 509176 421984 509182
rect 421932 509118 421984 509124
rect 421840 508836 421892 508842
rect 421840 508778 421892 508784
rect 421748 508768 421800 508774
rect 421748 508710 421800 508716
rect 421656 508700 421708 508706
rect 421656 508642 421708 508648
rect 414388 507884 414782 507890
rect 166814 507855 166870 507864
rect 414440 507878 414782 507884
rect 414388 507826 414440 507832
rect 236368 507816 236420 507822
rect 211554 507754 211936 507770
rect 227194 507754 227576 507770
rect 236118 507764 236368 507770
rect 236118 507758 236420 507764
rect 211554 507748 211948 507754
rect 211554 507742 211896 507748
rect 227194 507748 227588 507754
rect 227194 507742 227536 507748
rect 211896 507690 211948 507696
rect 236118 507742 236408 507758
rect 227536 507690 227588 507696
rect 218520 507680 218572 507686
rect 204838 507618 205128 507634
rect 209346 507618 209544 507634
rect 218270 507628 218520 507634
rect 218270 507622 218572 507628
rect 204838 507612 205140 507618
rect 204838 507606 205088 507612
rect 209346 507612 209556 507618
rect 209346 507606 209504 507612
rect 205088 507554 205140 507560
rect 218270 507606 218560 507622
rect 209504 507554 209556 507560
rect 202788 507544 202840 507550
rect 195808 507482 195914 507498
rect 195796 507476 195914 507482
rect 195848 507470 195914 507476
rect 202630 507492 202788 507498
rect 202630 507486 202840 507492
rect 202630 507470 202828 507486
rect 195796 507418 195848 507424
rect 191656 507408 191708 507414
rect 171598 507376 171654 507385
rect 171350 507334 171598 507362
rect 178406 507376 178462 507385
rect 178066 507334 178406 507362
rect 171598 507311 171654 507320
rect 182482 507346 182864 507362
rect 189198 507346 189488 507362
rect 191406 507356 191656 507362
rect 191406 507350 191708 507356
rect 182482 507340 182876 507346
rect 182482 507334 182824 507340
rect 178406 507311 178462 507320
rect 189198 507340 189500 507346
rect 189198 507334 189448 507340
rect 182824 507282 182876 507288
rect 191406 507334 191696 507350
rect 189448 507282 189500 507288
rect 184940 507272 184992 507278
rect 184782 507220 184940 507226
rect 184782 507214 184992 507220
rect 349712 507272 349764 507278
rect 349764 507220 350014 507226
rect 349712 507214 350014 507220
rect 184782 507198 184980 507214
rect 349724 507198 350014 507214
rect 421562 506560 421618 506569
rect 421562 506495 421618 506504
rect 165724 200926 166014 200954
rect 166184 200926 166474 200954
rect 167196 200926 167486 200954
rect 167656 200926 168038 200954
rect 168760 200926 169050 200954
rect 169312 200926 169602 200954
rect 169772 200926 170062 200954
rect 170232 200926 170614 200954
rect 171336 200926 171626 200954
rect 171704 200926 172178 200954
rect 172532 200926 172638 200954
rect 172808 200926 173190 200954
rect 173360 200926 173742 200954
rect 174004 200926 174202 200954
rect 174464 200926 174754 200954
rect 175476 200926 175766 200954
rect 175844 200926 176318 200954
rect 176948 200926 177330 200954
rect 177592 200926 177882 200954
rect 178052 200926 178342 200954
rect 178420 200926 178894 200954
rect 179064 200926 179354 200954
rect 179432 200926 179906 200954
rect 179984 200926 180458 200954
rect 180812 200926 180918 200954
rect 181088 200926 181470 200954
rect 181640 200926 181930 200954
rect 182192 200926 182482 200954
rect 182560 200926 183034 200954
rect 183112 200926 183494 200954
rect 183664 200926 184046 200954
rect 184216 200926 184598 200954
rect 185320 200926 185610 200954
rect 185688 200926 186070 200954
rect 186516 200926 186622 200954
rect 186792 200926 187174 200954
rect 187344 200926 187634 200954
rect 187712 200926 188186 200954
rect 188264 200926 188646 200954
rect 189092 200926 189198 200954
rect 189276 200926 189750 200954
rect 189920 200926 190210 200954
rect 190472 200926 190762 200954
rect 190840 200926 191314 200954
rect 191392 200926 191774 200954
rect 191944 200926 192326 200954
rect 192404 200926 192786 200954
rect 193600 200926 193890 200954
rect 193968 200926 194350 200954
rect 194704 200926 194902 200954
rect 195072 200926 195362 200954
rect 195440 200926 195914 200954
rect 196084 200926 196466 200954
rect 196544 200926 196926 200954
rect 197648 200926 197938 200954
rect 198200 200926 198490 200954
rect 198936 200926 199042 200954
rect 199120 200926 199502 200954
rect 199672 200926 200054 200954
rect 200132 200926 200606 200954
rect 200684 200926 201066 200954
rect 201512 200926 201618 200954
rect 201696 200926 202078 200954
rect 202248 200926 202630 200954
rect 202984 200926 203182 200954
rect 203352 200926 203642 200954
rect 203904 200926 204194 200954
rect 204272 200926 204654 200954
rect 204732 200926 205206 200954
rect 205652 200926 205758 200954
rect 205928 200926 206218 200954
rect 206388 200926 206770 200954
rect 207032 200926 207322 200954
rect 207400 200926 207782 200954
rect 207860 200926 208334 200954
rect 208504 200926 208794 200954
rect 208964 200926 209346 200954
rect 210068 200926 210358 200954
rect 210528 200926 210910 200954
rect 211632 200926 211922 200954
rect 212184 200926 212474 200954
rect 212644 200926 212934 200954
rect 213104 200926 213486 200954
rect 214116 200926 214498 200954
rect 214760 200926 215050 200954
rect 215312 200926 215510 200954
rect 215588 200926 216062 200954
rect 216232 200926 216614 200954
rect 216784 200926 217074 200954
rect 217152 200926 217626 200954
rect 218256 200926 218638 200954
rect 218716 200926 219190 200954
rect 219452 200926 219650 200954
rect 219912 200926 220202 200954
rect 220280 200926 220662 200954
rect 220832 200926 221214 200954
rect 221292 200926 221766 200954
rect 222396 200926 222778 200954
rect 222856 200926 223238 200954
rect 223684 200926 223790 200954
rect 223960 200926 224342 200954
rect 224512 200926 224802 200954
rect 225064 200926 225354 200954
rect 225432 200926 225906 200954
rect 226536 200926 226918 200954
rect 226996 200926 227378 200954
rect 227732 200926 227930 200954
rect 228008 200926 228482 200954
rect 228560 200926 228942 200954
rect 229204 200926 229494 200954
rect 229664 200926 229954 200954
rect 230676 200926 231058 200954
rect 231136 200926 231518 200954
rect 231964 200926 232070 200954
rect 232148 200926 232622 200954
rect 232792 200926 233082 200954
rect 233252 200926 233634 200954
rect 233712 200926 234094 200954
rect 234816 200926 235198 200954
rect 235276 200926 235658 200954
rect 236012 200926 236210 200954
rect 236288 200926 236670 200954
rect 236748 200926 237222 200954
rect 237484 200926 237774 200954
rect 237944 200926 238234 200954
rect 238956 200926 239246 200954
rect 239416 200926 239798 200954
rect 240520 200926 240810 200954
rect 241072 200926 241362 200954
rect 241532 200926 241914 200954
rect 241992 200926 242374 200954
rect 243096 200926 243386 200954
rect 243648 200926 243938 200954
rect 244660 200926 244950 200954
rect 245120 200926 245502 200954
rect 245856 200926 245962 200954
rect 246224 200926 246514 200954
rect 247236 200926 247526 200954
rect 247696 200926 248078 200954
rect 248432 200926 248630 200954
rect 248708 200926 249090 200954
rect 249168 200926 249642 200954
rect 249812 200926 250102 200954
rect 250180 200926 250654 200954
rect 251468 200926 251666 200954
rect 251928 200926 252218 200954
rect 252848 200926 253230 200954
rect 253308 200926 253782 200954
rect 253952 200926 254242 200954
rect 254320 200926 254794 200954
rect 254872 200926 255254 200954
rect 255424 200926 255806 200954
rect 255884 200926 256358 200954
rect 257080 200926 257370 200954
rect 257448 200926 257922 200954
rect 258184 200926 258382 200954
rect 258552 200926 258934 200954
rect 259012 200926 259394 200954
rect 259656 200926 259946 200954
rect 260208 200926 260498 200954
rect 261128 200926 261510 200954
rect 261680 200926 261970 200954
rect 262416 200926 262522 200954
rect 262784 200926 263074 200954
rect 263152 200926 263534 200954
rect 263704 200926 264086 200954
rect 264348 200926 264638 200954
rect 264992 200926 265098 200954
rect 265176 200926 265650 200954
rect 265728 200926 266110 200954
rect 266372 200926 266662 200954
rect 266740 200926 267214 200954
rect 267384 200926 267674 200954
rect 267936 200926 268226 200954
rect 268304 200926 268686 200954
rect 269132 200926 269238 200954
rect 269408 200926 269790 200954
rect 269960 200926 270250 200954
rect 270604 200926 270802 200954
rect 270880 200926 271262 200954
rect 271432 200926 271814 200954
rect 271984 200926 272366 200954
rect 272536 200926 272826 200954
rect 273640 200926 273930 200954
rect 274008 200926 274390 200954
rect 274836 200926 274942 200954
rect 275112 200926 275402 200954
rect 275664 200926 275954 200954
rect 276216 200926 276506 200954
rect 276584 200926 276966 200954
rect 277688 200926 277978 200954
rect 278240 200926 278530 200954
rect 278792 200926 279082 200954
rect 279160 200926 279542 200954
rect 279712 200926 280094 200954
rect 280356 200926 280554 200954
rect 280816 200926 281106 200954
rect 281552 200926 281658 200954
rect 281736 200926 282118 200954
rect 282288 200926 282670 200954
rect 282932 200926 283222 200954
rect 283392 200926 283682 200954
rect 283944 200926 284234 200954
rect 284312 200926 284694 200954
rect 284864 200926 285246 200954
rect 285692 200926 285798 200954
rect 285968 200926 286258 200954
rect 286520 200926 286810 200954
rect 287072 200926 287270 200954
rect 287440 200926 287822 200954
rect 287900 200926 288374 200954
rect 288544 200926 288834 200954
rect 289096 200926 289386 200954
rect 289832 200926 289938 200954
rect 290108 200926 290398 200954
rect 290568 200926 290950 200954
rect 291304 200926 291410 200954
rect 291672 200926 291962 200954
rect 292132 200926 292514 200954
rect 292592 200926 292974 200954
rect 293052 200926 293526 200954
rect 294248 200926 294538 200954
rect 321296 200926 321402 200954
rect 335096 200926 335294 200954
rect 339328 200926 339434 200954
rect 343376 200926 343574 200954
rect 347608 200926 347714 200954
rect 351748 200926 351854 200954
rect 355888 200926 355994 200954
rect 360028 200926 360134 200954
rect 364168 200926 364274 200954
rect 368308 200926 368414 200954
rect 372448 200926 372554 200954
rect 411088 200926 411194 200954
rect 415228 200926 415334 200954
rect 419368 200926 419474 200954
rect 101588 197872 101640 197878
rect 101588 197814 101640 197820
rect 101496 97980 101548 97986
rect 101496 97922 101548 97928
rect 101404 20664 101456 20670
rect 101404 20606 101456 20612
rect 101036 8152 101088 8158
rect 101036 8094 101088 8100
rect 98644 3732 98696 3738
rect 98644 3674 98696 3680
rect 99288 3732 99340 3738
rect 99288 3674 99340 3680
rect 99840 3732 99892 3738
rect 99840 3674 99892 3680
rect 98552 3120 98604 3126
rect 98552 3062 98604 3068
rect 98656 480 98684 3674
rect 99852 480 99880 3674
rect 101048 480 101076 8094
rect 101600 3738 101628 197814
rect 107568 197804 107620 197810
rect 107568 197746 107620 197752
rect 105544 197600 105596 197606
rect 105544 197542 105596 197548
rect 103428 89208 103480 89214
rect 103428 89150 103480 89156
rect 103440 3738 103468 89150
rect 104532 8220 104584 8226
rect 104532 8162 104584 8168
rect 101588 3732 101640 3738
rect 101588 3674 101640 3680
rect 102232 3732 102284 3738
rect 102232 3674 102284 3680
rect 103428 3732 103480 3738
rect 103428 3674 103480 3680
rect 102244 480 102272 3674
rect 103336 3120 103388 3126
rect 103336 3062 103388 3068
rect 103348 480 103376 3062
rect 104544 480 104572 8162
rect 105556 3058 105584 197542
rect 106188 86284 106240 86290
rect 106188 86226 106240 86232
rect 106200 3738 106228 86226
rect 107580 3738 107608 197746
rect 114468 197736 114520 197742
rect 114468 197678 114520 197684
rect 111064 197464 111116 197470
rect 111064 197406 111116 197412
rect 110328 17332 110380 17338
rect 110328 17274 110380 17280
rect 108120 8288 108172 8294
rect 108120 8230 108172 8236
rect 105728 3732 105780 3738
rect 105728 3674 105780 3680
rect 106188 3732 106240 3738
rect 106188 3674 106240 3680
rect 106924 3732 106976 3738
rect 106924 3674 106976 3680
rect 107568 3732 107620 3738
rect 107568 3674 107620 3680
rect 105544 3052 105596 3058
rect 105544 2994 105596 3000
rect 105740 480 105768 3674
rect 106936 480 106964 3674
rect 108132 480 108160 8230
rect 110340 3738 110368 17274
rect 109316 3732 109368 3738
rect 109316 3674 109368 3680
rect 110328 3732 110380 3738
rect 110328 3674 110380 3680
rect 109328 480 109356 3674
rect 110512 3052 110564 3058
rect 110512 2994 110564 3000
rect 110524 480 110552 2994
rect 111076 2990 111104 197406
rect 113088 84992 113140 84998
rect 113088 84934 113140 84940
rect 111616 7540 111668 7546
rect 111616 7482 111668 7488
rect 111064 2984 111116 2990
rect 111064 2926 111116 2932
rect 111628 480 111656 7482
rect 113100 6914 113128 84934
rect 112824 6886 113128 6914
rect 112824 480 112852 6886
rect 114480 3738 114508 197678
rect 125508 197532 125560 197538
rect 125508 197474 125560 197480
rect 124128 16244 124180 16250
rect 124128 16186 124180 16192
rect 119896 16176 119948 16182
rect 119896 16118 119948 16124
rect 117228 14748 117280 14754
rect 117228 14690 117280 14696
rect 115204 7472 115256 7478
rect 115204 7414 115256 7420
rect 114008 3732 114060 3738
rect 114008 3674 114060 3680
rect 114468 3732 114520 3738
rect 114468 3674 114520 3680
rect 114020 480 114048 3674
rect 115216 480 115244 7414
rect 117240 3738 117268 14690
rect 118792 7404 118844 7410
rect 118792 7346 118844 7352
rect 116400 3732 116452 3738
rect 116400 3674 116452 3680
rect 117228 3732 117280 3738
rect 117228 3674 117280 3680
rect 116412 480 116440 3674
rect 117596 2984 117648 2990
rect 117596 2926 117648 2932
rect 117608 480 117636 2926
rect 118804 480 118832 7346
rect 119908 480 119936 16118
rect 122288 7336 122340 7342
rect 122288 7278 122340 7284
rect 121092 2916 121144 2922
rect 121092 2858 121144 2864
rect 121104 480 121132 2858
rect 122300 480 122328 7278
rect 124140 3738 124168 16186
rect 125520 3738 125548 197474
rect 165620 195288 165672 195294
rect 165620 195230 165672 195236
rect 135168 87780 135220 87786
rect 135168 87722 135220 87728
rect 129648 17400 129700 17406
rect 129648 17342 129700 17348
rect 126888 14612 126940 14618
rect 126888 14554 126940 14560
rect 126900 3738 126928 14554
rect 129660 6914 129688 17342
rect 133788 17264 133840 17270
rect 133788 17206 133840 17212
rect 131028 13116 131080 13122
rect 131028 13058 131080 13064
rect 129384 6886 129688 6914
rect 128176 6112 128228 6118
rect 128176 6054 128228 6060
rect 126980 4480 127032 4486
rect 126980 4422 127032 4428
rect 123484 3732 123536 3738
rect 123484 3674 123536 3680
rect 124128 3732 124180 3738
rect 124128 3674 124180 3680
rect 124680 3732 124732 3738
rect 124680 3674 124732 3680
rect 125508 3732 125560 3738
rect 125508 3674 125560 3680
rect 125876 3732 125928 3738
rect 125876 3674 125928 3680
rect 126888 3732 126940 3738
rect 126888 3674 126940 3680
rect 123496 480 123524 3674
rect 124692 480 124720 3674
rect 125888 480 125916 3674
rect 126992 480 127020 4422
rect 128188 480 128216 6054
rect 129384 480 129412 6886
rect 131040 3738 131068 13058
rect 131764 9308 131816 9314
rect 131764 9250 131816 9256
rect 130568 3732 130620 3738
rect 130568 3674 130620 3680
rect 131028 3732 131080 3738
rect 131028 3674 131080 3680
rect 130580 480 130608 3674
rect 131776 480 131804 9250
rect 133800 3738 133828 17206
rect 135180 3738 135208 87722
rect 162768 85128 162820 85134
rect 162768 85070 162820 85076
rect 143448 85060 143500 85066
rect 143448 85002 143500 85008
rect 137928 84924 137980 84930
rect 137928 84866 137980 84872
rect 136456 9444 136508 9450
rect 136456 9386 136508 9392
rect 135260 9376 135312 9382
rect 135260 9318 135312 9324
rect 132960 3732 133012 3738
rect 132960 3674 133012 3680
rect 133788 3732 133840 3738
rect 133788 3674 133840 3680
rect 134156 3732 134208 3738
rect 134156 3674 134208 3680
rect 135168 3732 135220 3738
rect 135168 3674 135220 3680
rect 132972 480 133000 3674
rect 134168 480 134196 3674
rect 135272 480 135300 9318
rect 136468 480 136496 9386
rect 137940 6914 137968 84866
rect 140688 18624 140740 18630
rect 140688 18566 140740 18572
rect 139308 16040 139360 16046
rect 139308 15982 139360 15988
rect 137664 6886 137968 6914
rect 137664 480 137692 6886
rect 139320 3738 139348 15982
rect 140700 3738 140728 18566
rect 141240 6044 141292 6050
rect 141240 5986 141292 5992
rect 138848 3732 138900 3738
rect 138848 3674 138900 3680
rect 139308 3732 139360 3738
rect 139308 3674 139360 3680
rect 140044 3732 140096 3738
rect 140044 3674 140096 3680
rect 140688 3732 140740 3738
rect 140688 3674 140740 3680
rect 138860 480 138888 3674
rect 140056 480 140084 3674
rect 141252 480 141280 5986
rect 143460 3738 143488 85002
rect 147588 80708 147640 80714
rect 147588 80650 147640 80656
rect 144828 17468 144880 17474
rect 144828 17410 144880 17416
rect 144736 5976 144788 5982
rect 144736 5918 144788 5924
rect 142436 3732 142488 3738
rect 142436 3674 142488 3680
rect 143448 3732 143500 3738
rect 143448 3674 143500 3680
rect 143540 3732 143592 3738
rect 143540 3674 143592 3680
rect 142448 480 142476 3674
rect 143552 480 143580 3674
rect 144748 480 144776 5918
rect 144840 3738 144868 17410
rect 145932 13184 145984 13190
rect 145932 13126 145984 13132
rect 144828 3732 144880 3738
rect 144828 3674 144880 3680
rect 145944 480 145972 13126
rect 147600 3738 147628 80650
rect 161388 17536 161440 17542
rect 161388 17478 161440 17484
rect 149520 7268 149572 7274
rect 149520 7210 149572 7216
rect 148324 5908 148376 5914
rect 148324 5850 148376 5856
rect 147128 3732 147180 3738
rect 147128 3674 147180 3680
rect 147588 3732 147640 3738
rect 147588 3674 147640 3680
rect 147140 480 147168 3674
rect 148336 480 148364 5850
rect 149532 480 149560 7210
rect 153016 7200 153068 7206
rect 153016 7142 153068 7148
rect 151820 5840 151872 5846
rect 151820 5782 151872 5788
rect 150624 4412 150676 4418
rect 150624 4354 150676 4360
rect 150636 480 150664 4354
rect 151832 480 151860 5782
rect 153028 480 153056 7142
rect 156604 7132 156656 7138
rect 156604 7074 156656 7080
rect 155408 5772 155460 5778
rect 155408 5714 155460 5720
rect 154212 4344 154264 4350
rect 154212 4286 154264 4292
rect 154224 480 154252 4286
rect 155420 480 155448 5714
rect 156616 480 156644 7074
rect 160100 7064 160152 7070
rect 160100 7006 160152 7012
rect 158904 5704 158956 5710
rect 158904 5646 158956 5652
rect 157800 4276 157852 4282
rect 157800 4218 157852 4224
rect 157812 480 157840 4218
rect 158916 480 158944 5646
rect 160112 480 160140 7006
rect 161400 6914 161428 17478
rect 162780 6914 162808 85070
rect 165528 16108 165580 16114
rect 165528 16050 165580 16056
rect 161308 6886 161428 6914
rect 162504 6886 162808 6914
rect 161308 480 161336 6886
rect 162504 480 162532 6886
rect 163688 5636 163740 5642
rect 163688 5578 163740 5584
rect 163700 480 163728 5578
rect 165540 3466 165568 16050
rect 165632 4894 165660 195230
rect 165620 4888 165672 4894
rect 165620 4830 165672 4836
rect 165724 4826 165752 200926
rect 166184 195294 166212 200926
rect 167026 200790 167132 200818
rect 167104 200114 167132 200790
rect 167012 200086 167132 200114
rect 166172 195288 166224 195294
rect 166172 195230 166224 195236
rect 166908 14680 166960 14686
rect 166908 14622 166960 14628
rect 165712 4820 165764 4826
rect 165712 4762 165764 4768
rect 166920 3466 166948 14622
rect 167012 4962 167040 200086
rect 167196 180794 167224 200926
rect 167656 198082 167684 200926
rect 168590 200790 168696 200818
rect 168472 200456 168524 200462
rect 168472 200398 168524 200404
rect 167644 198076 167696 198082
rect 167644 198018 167696 198024
rect 168380 192024 168432 192030
rect 168380 191966 168432 191972
rect 167104 180766 167224 180794
rect 167104 6186 167132 180766
rect 168392 6254 168420 191966
rect 168380 6248 168432 6254
rect 168380 6190 168432 6196
rect 167092 6180 167144 6186
rect 167092 6122 167144 6128
rect 167184 6180 167236 6186
rect 167184 6122 167236 6128
rect 167000 4956 167052 4962
rect 167000 4898 167052 4904
rect 164884 3460 164936 3466
rect 164884 3402 164936 3408
rect 165528 3460 165580 3466
rect 165528 3402 165580 3408
rect 166080 3460 166132 3466
rect 166080 3402 166132 3408
rect 166908 3460 166960 3466
rect 166908 3402 166960 3408
rect 164896 480 164924 3402
rect 166092 480 166120 3402
rect 167196 480 167224 6122
rect 168484 5030 168512 200398
rect 168472 5024 168524 5030
rect 168472 4966 168524 4972
rect 168668 3738 168696 200790
rect 168760 200462 168788 200926
rect 168748 200456 168800 200462
rect 168748 200398 168800 200404
rect 169312 192030 169340 200926
rect 169772 198014 169800 200926
rect 170232 198150 170260 200926
rect 171166 200790 171272 200818
rect 170220 198144 170272 198150
rect 170220 198086 170272 198092
rect 169760 198008 169812 198014
rect 169760 197950 169812 197956
rect 170404 198008 170456 198014
rect 170404 197950 170456 197956
rect 169576 196852 169628 196858
rect 169576 196794 169628 196800
rect 169300 192024 169352 192030
rect 169300 191966 169352 191972
rect 168656 3732 168708 3738
rect 168656 3674 168708 3680
rect 169588 3466 169616 196794
rect 170416 89078 170444 197950
rect 170404 89072 170456 89078
rect 170404 89014 170456 89020
rect 170772 6248 170824 6254
rect 170772 6190 170824 6196
rect 169668 5160 169720 5166
rect 169668 5102 169720 5108
rect 168380 3460 168432 3466
rect 168380 3402 168432 3408
rect 169576 3460 169628 3466
rect 169576 3402 169628 3408
rect 168392 480 168420 3402
rect 169680 2666 169708 5102
rect 169588 2638 169708 2666
rect 169588 480 169616 2638
rect 170784 480 170812 6190
rect 171244 5098 171272 200790
rect 171336 196654 171364 200926
rect 171324 196648 171376 196654
rect 171324 196590 171376 196596
rect 171704 180794 171732 200926
rect 171336 180766 171732 180794
rect 171232 5092 171284 5098
rect 171232 5034 171284 5040
rect 171336 3534 171364 180766
rect 171968 9512 172020 9518
rect 171968 9454 172020 9460
rect 171324 3528 171376 3534
rect 171324 3470 171376 3476
rect 171980 480 172008 9454
rect 172532 3602 172560 200926
rect 172704 195288 172756 195294
rect 172704 195230 172756 195236
rect 172716 14482 172744 195230
rect 172704 14476 172756 14482
rect 172704 14418 172756 14424
rect 172808 4214 172836 200926
rect 173164 197396 173216 197402
rect 173164 197338 173216 197344
rect 173176 87650 173204 197338
rect 173360 195294 173388 200926
rect 174004 198218 174032 200926
rect 174464 198694 174492 200926
rect 175306 200790 175412 200818
rect 174452 198688 174504 198694
rect 174452 198630 174504 198636
rect 173992 198212 174044 198218
rect 173992 198154 174044 198160
rect 173348 195288 173400 195294
rect 173348 195230 173400 195236
rect 173164 87644 173216 87650
rect 173164 87586 173216 87592
rect 175384 6322 175412 200790
rect 175476 89010 175504 200926
rect 175844 180794 175872 200926
rect 176778 200790 176884 200818
rect 175568 180766 175872 180794
rect 175464 89004 175516 89010
rect 175464 88946 175516 88952
rect 175464 9580 175516 9586
rect 175464 9522 175516 9528
rect 175372 6316 175424 6322
rect 175372 6258 175424 6264
rect 173164 5092 173216 5098
rect 173164 5034 173216 5040
rect 172796 4208 172848 4214
rect 172796 4150 172848 4156
rect 172520 3596 172572 3602
rect 172520 3538 172572 3544
rect 173176 480 173204 5034
rect 174268 4820 174320 4826
rect 174268 4762 174320 4768
rect 174280 480 174308 4762
rect 175476 480 175504 9522
rect 175568 3670 175596 180766
rect 176660 3732 176712 3738
rect 176660 3674 176712 3680
rect 175556 3664 175608 3670
rect 175556 3606 175608 3612
rect 176672 480 176700 3674
rect 176856 2854 176884 200790
rect 176948 6390 176976 200926
rect 177304 198688 177356 198694
rect 177304 198630 177356 198636
rect 177316 16182 177344 198630
rect 177592 197402 177620 200926
rect 178052 198286 178080 200926
rect 178040 198280 178092 198286
rect 178040 198222 178092 198228
rect 177580 197396 177632 197402
rect 177580 197338 177632 197344
rect 178132 195288 178184 195294
rect 178132 195230 178184 195236
rect 178144 22778 178172 195230
rect 178420 180794 178448 200926
rect 178684 198280 178736 198286
rect 178684 198222 178736 198228
rect 178236 180766 178448 180794
rect 178132 22772 178184 22778
rect 178132 22714 178184 22720
rect 177304 16176 177356 16182
rect 177304 16118 177356 16124
rect 178236 6458 178264 180766
rect 178696 16250 178724 198222
rect 179064 195294 179092 200926
rect 179052 195288 179104 195294
rect 179052 195230 179104 195236
rect 178684 16244 178736 16250
rect 178684 16186 178736 16192
rect 178224 6452 178276 6458
rect 178224 6394 178276 6400
rect 176936 6384 176988 6390
rect 176936 6326 176988 6332
rect 177856 4208 177908 4214
rect 177856 4150 177908 4156
rect 176844 2848 176896 2854
rect 176844 2790 176896 2796
rect 177868 480 177896 4150
rect 179432 3670 179460 200926
rect 179984 180794 180012 200926
rect 180812 198014 180840 200926
rect 181088 198422 181116 200926
rect 181640 200114 181668 200926
rect 181272 200086 181668 200114
rect 181076 198416 181128 198422
rect 181076 198358 181128 198364
rect 180800 198008 180852 198014
rect 180800 197950 180852 197956
rect 180064 196648 180116 196654
rect 180064 196590 180116 196596
rect 179524 180766 180012 180794
rect 179524 6526 179552 180766
rect 179512 6520 179564 6526
rect 179512 6462 179564 6468
rect 179420 3664 179472 3670
rect 179420 3606 179472 3612
rect 180076 3534 180104 196590
rect 181272 180794 181300 200086
rect 181444 197396 181496 197402
rect 181444 197338 181496 197344
rect 180996 180766 181300 180794
rect 180996 6594 181024 180766
rect 181456 15910 181484 197338
rect 182192 196722 182220 200926
rect 182180 196716 182232 196722
rect 182180 196658 182232 196664
rect 182272 195288 182324 195294
rect 182272 195230 182324 195236
rect 181444 15904 181496 15910
rect 181444 15846 181496 15852
rect 182284 6662 182312 195230
rect 182560 180794 182588 200926
rect 182824 198008 182876 198014
rect 182824 197950 182876 197956
rect 182376 180766 182588 180794
rect 182272 6656 182324 6662
rect 182272 6598 182324 6604
rect 180984 6588 181036 6594
rect 180984 6530 181036 6536
rect 182376 3806 182404 180766
rect 182836 3874 182864 197950
rect 183112 195294 183140 200926
rect 183100 195288 183152 195294
rect 183100 195230 183152 195236
rect 183664 87718 183692 200926
rect 184216 198490 184244 200926
rect 185058 200790 185164 200818
rect 184204 198484 184256 198490
rect 184204 198426 184256 198432
rect 184296 198484 184348 198490
rect 184296 198426 184348 198432
rect 184204 198076 184256 198082
rect 184204 198018 184256 198024
rect 183652 87712 183704 87718
rect 183652 87654 183704 87660
rect 184216 4078 184244 198018
rect 184308 4146 184336 198426
rect 184388 198212 184440 198218
rect 184388 198154 184440 198160
rect 184400 14754 184428 198154
rect 185136 180794 185164 200790
rect 185320 197402 185348 200926
rect 185688 200114 185716 200926
rect 185504 200086 185716 200114
rect 185308 197396 185360 197402
rect 185308 197338 185360 197344
rect 185504 180794 185532 200086
rect 185584 198416 185636 198422
rect 185584 198358 185636 198364
rect 185044 180766 185164 180794
rect 185228 180766 185532 180794
rect 184388 14748 184440 14754
rect 184388 14690 184440 14696
rect 185044 6730 185072 180766
rect 185032 6724 185084 6730
rect 185032 6666 185084 6672
rect 184296 4140 184348 4146
rect 184296 4082 184348 4088
rect 184204 4072 184256 4078
rect 184204 4014 184256 4020
rect 185228 4010 185256 180766
rect 185216 4004 185268 4010
rect 185216 3946 185268 3952
rect 182824 3868 182876 3874
rect 182824 3810 182876 3816
rect 182364 3800 182416 3806
rect 182364 3742 182416 3748
rect 184940 3800 184992 3806
rect 184940 3742 184992 3748
rect 180248 3664 180300 3670
rect 180248 3606 180300 3612
rect 179052 3528 179104 3534
rect 179052 3470 179104 3476
rect 180064 3528 180116 3534
rect 180064 3470 180116 3476
rect 179064 480 179092 3470
rect 180260 480 180288 3606
rect 183744 3460 183796 3466
rect 183744 3402 183796 3408
rect 181444 3392 181496 3398
rect 181444 3334 181496 3340
rect 181456 480 181484 3334
rect 182548 2848 182600 2854
rect 182548 2790 182600 2796
rect 182560 480 182588 2790
rect 183756 480 183784 3402
rect 184952 480 184980 3742
rect 185596 3534 185624 198358
rect 186412 195288 186464 195294
rect 186412 195230 186464 195236
rect 186424 7614 186452 195230
rect 186412 7608 186464 7614
rect 186412 7550 186464 7556
rect 186516 5234 186544 200926
rect 186792 195294 186820 200926
rect 187344 198014 187372 200926
rect 187332 198008 187384 198014
rect 187332 197950 187384 197956
rect 186964 197396 187016 197402
rect 186964 197338 187016 197344
rect 186780 195288 186832 195294
rect 186780 195230 186832 195236
rect 186504 5228 186556 5234
rect 186504 5170 186556 5176
rect 185584 3528 185636 3534
rect 185584 3470 185636 3476
rect 186136 3528 186188 3534
rect 186136 3470 186188 3476
rect 186148 480 186176 3470
rect 186976 3330 187004 197338
rect 187332 6316 187384 6322
rect 187332 6258 187384 6264
rect 186964 3324 187016 3330
rect 186964 3266 187016 3272
rect 187344 480 187372 6258
rect 187712 5302 187740 200926
rect 188264 180794 188292 200926
rect 189092 198354 189120 200926
rect 189080 198348 189132 198354
rect 189080 198290 189132 198296
rect 188344 196716 188396 196722
rect 188344 196658 188396 196664
rect 187804 180766 188292 180794
rect 187804 7682 187832 180766
rect 187792 7676 187844 7682
rect 187792 7618 187844 7624
rect 187700 5296 187752 5302
rect 187700 5238 187752 5244
rect 188356 3534 188384 196658
rect 189276 5370 189304 200926
rect 189920 200114 189948 200926
rect 189368 200086 189948 200114
rect 189368 7750 189396 200086
rect 190472 198082 190500 200926
rect 190460 198076 190512 198082
rect 190460 198018 190512 198024
rect 189724 198008 189776 198014
rect 189724 197950 189776 197956
rect 189356 7744 189408 7750
rect 189356 7686 189408 7692
rect 189736 6914 189764 197950
rect 190552 195084 190604 195090
rect 190552 195026 190604 195032
rect 190564 7818 190592 195026
rect 190840 180794 190868 200926
rect 191104 198144 191156 198150
rect 191104 198086 191156 198092
rect 190656 180766 190868 180794
rect 190552 7812 190604 7818
rect 190552 7754 190604 7760
rect 189644 6886 189764 6914
rect 189264 5364 189316 5370
rect 189264 5306 189316 5312
rect 188528 3596 188580 3602
rect 188528 3538 188580 3544
rect 188344 3528 188396 3534
rect 188344 3470 188396 3476
rect 188540 480 188568 3538
rect 189644 3262 189672 6886
rect 190656 5438 190684 180766
rect 190828 6384 190880 6390
rect 190828 6326 190880 6332
rect 190644 5432 190696 5438
rect 190644 5374 190696 5380
rect 189724 4888 189776 4894
rect 189724 4830 189776 4836
rect 189632 3256 189684 3262
rect 189632 3198 189684 3204
rect 189736 480 189764 4830
rect 190840 480 190868 6326
rect 191116 3194 191144 198086
rect 191392 195090 191420 200926
rect 191944 198558 191972 200926
rect 191932 198552 191984 198558
rect 191932 198494 191984 198500
rect 191380 195084 191432 195090
rect 191380 195026 191432 195032
rect 192404 180794 192432 200926
rect 193338 200790 193444 200818
rect 193416 200114 193444 200790
rect 193324 200086 193444 200114
rect 192484 198076 192536 198082
rect 192484 198018 192536 198024
rect 191944 180766 192432 180794
rect 191944 5506 191972 180766
rect 191932 5500 191984 5506
rect 191932 5442 191984 5448
rect 192024 3936 192076 3942
rect 192024 3878 192076 3884
rect 191104 3188 191156 3194
rect 191104 3130 191156 3136
rect 192036 480 192064 3878
rect 192496 3126 192524 198018
rect 193324 8974 193352 200086
rect 193600 198490 193628 200926
rect 193968 200114 193996 200926
rect 193784 200086 193996 200114
rect 193588 198484 193640 198490
rect 193588 198426 193640 198432
rect 193784 180794 193812 200086
rect 193864 198348 193916 198354
rect 193864 198290 193916 198296
rect 193416 180766 193812 180794
rect 193312 8968 193364 8974
rect 193312 8910 193364 8916
rect 193220 4956 193272 4962
rect 193220 4898 193272 4904
rect 192484 3120 192536 3126
rect 192484 3062 192536 3068
rect 193232 480 193260 4898
rect 193416 4758 193444 180766
rect 193404 4752 193456 4758
rect 193404 4694 193456 4700
rect 193876 3058 193904 198290
rect 194704 9042 194732 200926
rect 195072 198626 195100 200926
rect 195440 200114 195468 200926
rect 195164 200086 195468 200114
rect 195060 198620 195112 198626
rect 195060 198562 195112 198568
rect 195164 180794 195192 200086
rect 195244 198484 195296 198490
rect 195244 198426 195296 198432
rect 194796 180766 195192 180794
rect 194692 9036 194744 9042
rect 194692 8978 194744 8984
rect 194416 6452 194468 6458
rect 194416 6394 194468 6400
rect 193864 3052 193916 3058
rect 193864 2994 193916 3000
rect 194428 480 194456 6394
rect 194796 4622 194824 180766
rect 194784 4616 194836 4622
rect 194784 4558 194836 4564
rect 195256 2990 195284 198426
rect 196084 9110 196112 200926
rect 196544 198422 196572 200926
rect 197478 200790 197584 200818
rect 196900 198620 196952 198626
rect 196900 198562 196952 198568
rect 196532 198416 196584 198422
rect 196532 198358 196584 198364
rect 196808 198348 196860 198354
rect 196808 198290 196860 198296
rect 196820 195974 196848 198290
rect 196636 195946 196848 195974
rect 196072 9104 196124 9110
rect 196072 9046 196124 9052
rect 195244 2984 195296 2990
rect 195244 2926 195296 2932
rect 195612 2984 195664 2990
rect 195612 2926 195664 2932
rect 195624 480 195652 2926
rect 196636 2922 196664 195946
rect 196912 186314 196940 198562
rect 196728 186286 196940 186314
rect 196728 17338 196756 186286
rect 196716 17332 196768 17338
rect 196716 17274 196768 17280
rect 196808 17332 196860 17338
rect 196808 17274 196860 17280
rect 196820 6914 196848 17274
rect 196728 6886 196848 6914
rect 196624 2916 196676 2922
rect 196624 2858 196676 2864
rect 196728 2854 196756 6886
rect 196808 5024 196860 5030
rect 196808 4966 196860 4972
rect 196716 2848 196768 2854
rect 196716 2790 196768 2796
rect 196820 480 196848 4966
rect 197556 4690 197584 200790
rect 197648 9178 197676 200926
rect 198004 198552 198056 198558
rect 198004 198494 198056 198500
rect 198016 84998 198044 198494
rect 198200 197674 198228 200926
rect 198188 197668 198240 197674
rect 198188 197610 198240 197616
rect 198936 191282 198964 200926
rect 199120 200114 199148 200926
rect 199028 200086 199148 200114
rect 198924 191276 198976 191282
rect 198924 191218 198976 191224
rect 198924 191072 198976 191078
rect 198924 191014 198976 191020
rect 198832 188420 198884 188426
rect 198832 188362 198884 188368
rect 198004 84992 198056 84998
rect 198004 84934 198056 84940
rect 198096 84992 198148 84998
rect 198096 84934 198148 84940
rect 197636 9172 197688 9178
rect 197636 9114 197688 9120
rect 197912 6520 197964 6526
rect 197912 6462 197964 6468
rect 197544 4684 197596 4690
rect 197544 4626 197596 4632
rect 197924 480 197952 6462
rect 198108 2990 198136 84934
rect 198844 9246 198872 188362
rect 198832 9240 198884 9246
rect 198832 9182 198884 9188
rect 198936 4554 198964 191014
rect 199028 188426 199056 200086
rect 199384 197668 199436 197674
rect 199384 197610 199436 197616
rect 199016 188420 199068 188426
rect 199016 188362 199068 188368
rect 199396 86290 199424 197610
rect 199672 197402 199700 200926
rect 199660 197396 199712 197402
rect 199660 197338 199712 197344
rect 199384 86284 199436 86290
rect 199384 86226 199436 86232
rect 200132 6798 200160 200926
rect 200684 180794 200712 200926
rect 201512 197606 201540 200926
rect 201500 197600 201552 197606
rect 201500 197542 201552 197548
rect 200764 196920 200816 196926
rect 200764 196862 200816 196868
rect 200224 180766 200712 180794
rect 200224 89146 200252 180766
rect 200212 89140 200264 89146
rect 200212 89082 200264 89088
rect 200120 6792 200172 6798
rect 200120 6734 200172 6740
rect 200304 4752 200356 4758
rect 200304 4694 200356 4700
rect 198924 4548 198976 4554
rect 198924 4490 198976 4496
rect 199108 3868 199160 3874
rect 199108 3810 199160 3816
rect 198096 2984 198148 2990
rect 198096 2926 198148 2932
rect 199120 480 199148 3810
rect 200316 480 200344 4694
rect 200776 3738 200804 196862
rect 201696 6866 201724 200926
rect 202248 200114 202276 200926
rect 201788 200086 202276 200114
rect 201788 14550 201816 200086
rect 202144 197464 202196 197470
rect 202144 197406 202196 197412
rect 202156 44878 202184 197406
rect 202984 197402 203012 200926
rect 202972 197396 203024 197402
rect 202972 197338 203024 197344
rect 203352 180794 203380 200926
rect 203904 196790 203932 200926
rect 204272 198014 204300 200926
rect 204260 198008 204312 198014
rect 204260 197950 204312 197956
rect 203892 196784 203944 196790
rect 203892 196726 203944 196732
rect 204732 180794 204760 200926
rect 205652 197402 205680 200926
rect 205928 197946 205956 200926
rect 206388 200114 206416 200926
rect 206204 200086 206416 200114
rect 205916 197940 205968 197946
rect 205916 197882 205968 197888
rect 204904 197396 204956 197402
rect 204904 197338 204956 197344
rect 205640 197396 205692 197402
rect 205640 197338 205692 197344
rect 203076 180766 203380 180794
rect 204364 180766 204760 180794
rect 202144 44872 202196 44878
rect 202144 44814 202196 44820
rect 202788 22772 202840 22778
rect 202788 22714 202840 22720
rect 201776 14544 201828 14550
rect 201776 14486 201828 14492
rect 202144 14476 202196 14482
rect 202144 14418 202196 14424
rect 201684 6860 201736 6866
rect 201684 6802 201736 6808
rect 201500 6588 201552 6594
rect 201500 6530 201552 6536
rect 200764 3732 200816 3738
rect 200764 3674 200816 3680
rect 201512 480 201540 6530
rect 202156 3806 202184 14418
rect 202800 6914 202828 22714
rect 203076 7886 203104 180766
rect 204364 7954 204392 180766
rect 204916 15978 204944 197338
rect 206204 180794 206232 200086
rect 206928 198008 206980 198014
rect 206928 197950 206980 197956
rect 206284 197396 206336 197402
rect 206284 197338 206336 197344
rect 205836 180766 206232 180794
rect 204996 155236 205048 155242
rect 204996 155178 205048 155184
rect 204904 15972 204956 15978
rect 204904 15914 204956 15920
rect 204352 7948 204404 7954
rect 204352 7890 204404 7896
rect 203064 7880 203116 7886
rect 203064 7822 203116 7828
rect 205008 6914 205036 155178
rect 205088 15904 205140 15910
rect 205088 15846 205140 15852
rect 202708 6886 202828 6914
rect 204916 6886 205036 6914
rect 202144 3800 202196 3806
rect 202144 3742 202196 3748
rect 202708 480 202736 6886
rect 203892 4684 203944 4690
rect 203892 4626 203944 4632
rect 203904 480 203932 4626
rect 204916 3670 204944 6886
rect 205100 3942 205128 15846
rect 205836 8022 205864 180766
rect 206296 84862 206324 197338
rect 206376 86284 206428 86290
rect 206376 86226 206428 86232
rect 206284 84856 206336 84862
rect 206284 84798 206336 84804
rect 205824 8016 205876 8022
rect 205824 7958 205876 7964
rect 205180 6656 205232 6662
rect 205180 6598 205232 6604
rect 205088 3936 205140 3942
rect 205088 3878 205140 3884
rect 204904 3664 204956 3670
rect 204904 3606 204956 3612
rect 205192 3346 205220 6598
rect 206388 3874 206416 86226
rect 206376 3868 206428 3874
rect 206376 3810 206428 3816
rect 206940 3398 206968 197950
rect 207032 197402 207060 200926
rect 207400 198150 207428 200926
rect 207388 198144 207440 198150
rect 207388 198086 207440 198092
rect 207020 197396 207072 197402
rect 207020 197338 207072 197344
rect 207860 180794 207888 200926
rect 208504 197470 208532 200926
rect 208964 197878 208992 200926
rect 209898 200790 210004 200818
rect 209044 197940 209096 197946
rect 209044 197882 209096 197888
rect 208952 197872 209004 197878
rect 208952 197814 209004 197820
rect 208492 197464 208544 197470
rect 208492 197406 208544 197412
rect 207216 180766 207888 180794
rect 207216 8090 207244 180766
rect 207204 8084 207256 8090
rect 207204 8026 207256 8032
rect 207388 5228 207440 5234
rect 207388 5170 207440 5176
rect 205100 3318 205220 3346
rect 206192 3392 206244 3398
rect 206192 3334 206244 3340
rect 206928 3392 206980 3398
rect 206928 3334 206980 3340
rect 205100 480 205128 3318
rect 206204 480 206232 3334
rect 207400 480 207428 5170
rect 209056 5098 209084 197882
rect 209136 197872 209188 197878
rect 209136 197814 209188 197820
rect 209148 5166 209176 197814
rect 209688 177336 209740 177342
rect 209688 177278 209740 177284
rect 209136 5160 209188 5166
rect 209136 5102 209188 5108
rect 209044 5092 209096 5098
rect 209044 5034 209096 5040
rect 209700 3398 209728 177278
rect 209976 8158 210004 200790
rect 210068 89214 210096 200926
rect 210528 198082 210556 200926
rect 211370 200790 211476 200818
rect 210516 198076 210568 198082
rect 210516 198018 210568 198024
rect 210976 198076 211028 198082
rect 210976 198018 211028 198024
rect 210056 89208 210108 89214
rect 210056 89150 210108 89156
rect 209964 8152 210016 8158
rect 209964 8094 210016 8100
rect 210988 3398 211016 198018
rect 211448 180794 211476 200790
rect 211632 197674 211660 200926
rect 212184 197810 212212 200926
rect 212172 197804 212224 197810
rect 212172 197746 212224 197752
rect 211620 197668 211672 197674
rect 211620 197610 211672 197616
rect 211356 180766 211476 180794
rect 211356 8226 211384 180766
rect 212644 8294 212672 200926
rect 213104 198626 213132 200926
rect 213946 200790 214052 200818
rect 213092 198620 213144 198626
rect 213092 198562 213144 198568
rect 213276 198620 213328 198626
rect 213276 198562 213328 198568
rect 213184 197668 213236 197674
rect 213184 197610 213236 197616
rect 213196 17542 213224 197610
rect 213288 80714 213316 198562
rect 214024 198490 214052 200790
rect 214012 198484 214064 198490
rect 214012 198426 214064 198432
rect 213828 198144 213880 198150
rect 213828 198086 213880 198092
rect 213276 80708 213328 80714
rect 213276 80650 213328 80656
rect 213184 17536 213236 17542
rect 213184 17478 213236 17484
rect 212632 8288 212684 8294
rect 212632 8230 212684 8236
rect 211344 8220 211396 8226
rect 211344 8162 211396 8168
rect 211068 5296 211120 5302
rect 211068 5238 211120 5244
rect 208584 3392 208636 3398
rect 208584 3334 208636 3340
rect 209688 3392 209740 3398
rect 209688 3334 209740 3340
rect 209780 3392 209832 3398
rect 209780 3334 209832 3340
rect 210976 3392 211028 3398
rect 210976 3334 211028 3340
rect 208596 480 208624 3334
rect 209792 480 209820 3334
rect 211080 2666 211108 5238
rect 212172 3664 212224 3670
rect 212172 3606 212224 3612
rect 210988 2638 211108 2666
rect 210988 480 211016 2638
rect 212184 480 212212 3606
rect 213840 3398 213868 198086
rect 214116 7546 214144 200926
rect 214760 198558 214788 200926
rect 214748 198552 214800 198558
rect 214748 198494 214800 198500
rect 214656 198484 214708 198490
rect 214656 198426 214708 198432
rect 214564 197804 214616 197810
rect 214564 197746 214616 197752
rect 214576 9450 214604 197746
rect 214668 18630 214696 198426
rect 215312 197742 215340 200926
rect 215300 197736 215352 197742
rect 215300 197678 215352 197684
rect 214656 18624 214708 18630
rect 214656 18566 214708 18572
rect 214564 9444 214616 9450
rect 214564 9386 214616 9392
rect 214104 7540 214156 7546
rect 214104 7482 214156 7488
rect 215588 7478 215616 200926
rect 216232 198218 216260 200926
rect 216784 198422 216812 200926
rect 216772 198416 216824 198422
rect 216772 198358 216824 198364
rect 216220 198212 216272 198218
rect 216220 198154 216272 198160
rect 216036 197736 216088 197742
rect 216036 197678 216088 197684
rect 215944 197600 215996 197606
rect 215944 197542 215996 197548
rect 215956 17406 215984 197542
rect 216048 85134 216076 197678
rect 217152 180794 217180 200926
rect 218086 200790 218192 200818
rect 218164 198694 218192 200790
rect 218152 198688 218204 198694
rect 218152 198630 218204 198636
rect 217324 198552 217376 198558
rect 217324 198494 217376 198500
rect 216784 180766 217180 180794
rect 216036 85128 216088 85134
rect 216036 85070 216088 85076
rect 216588 22840 216640 22846
rect 216588 22782 216640 22788
rect 215944 17400 215996 17406
rect 215944 17342 215996 17348
rect 215576 7472 215628 7478
rect 215576 7414 215628 7420
rect 214472 5364 214524 5370
rect 214472 5306 214524 5312
rect 213368 3392 213420 3398
rect 213368 3334 213420 3340
rect 213828 3392 213880 3398
rect 213828 3334 213880 3340
rect 213380 480 213408 3334
rect 214484 480 214512 5306
rect 216600 3398 216628 22782
rect 216784 7410 216812 180766
rect 217336 85066 217364 198494
rect 218256 198354 218284 200926
rect 218244 198348 218296 198354
rect 218244 198290 218296 198296
rect 217968 198212 218020 198218
rect 217968 198154 218020 198160
rect 217324 85060 217376 85066
rect 217324 85002 217376 85008
rect 216772 7404 216824 7410
rect 216772 7346 216824 7352
rect 217980 3398 218008 198154
rect 218716 180794 218744 200926
rect 219452 198286 219480 200926
rect 219440 198280 219492 198286
rect 219440 198222 219492 198228
rect 219912 197538 219940 200926
rect 220280 200114 220308 200926
rect 220096 200086 220308 200114
rect 219900 197532 219952 197538
rect 219900 197474 219952 197480
rect 220096 180794 220124 200086
rect 220728 198280 220780 198286
rect 220728 198222 220780 198228
rect 220176 197396 220228 197402
rect 220176 197338 220228 197344
rect 218256 180766 218744 180794
rect 219728 180766 220124 180794
rect 218256 7342 218284 180766
rect 219728 14618 219756 180766
rect 220084 171828 220136 171834
rect 220084 171770 220136 171776
rect 219716 14612 219768 14618
rect 219716 14554 219768 14560
rect 218244 7336 218296 7342
rect 218244 7278 218296 7284
rect 218060 5432 218112 5438
rect 218060 5374 218112 5380
rect 215668 3392 215720 3398
rect 215668 3334 215720 3340
rect 216588 3392 216640 3398
rect 216588 3334 216640 3340
rect 216864 3392 216916 3398
rect 216864 3334 216916 3340
rect 217968 3392 218020 3398
rect 217968 3334 218020 3340
rect 215680 480 215708 3334
rect 216876 480 216904 3334
rect 218072 480 218100 5374
rect 219256 3868 219308 3874
rect 219256 3810 219308 3816
rect 219268 480 219296 3810
rect 220096 3670 220124 171770
rect 220188 87786 220216 197338
rect 220176 87780 220228 87786
rect 220176 87722 220228 87728
rect 220740 6914 220768 198222
rect 220464 6886 220768 6914
rect 220084 3664 220136 3670
rect 220084 3606 220136 3612
rect 220464 480 220492 6886
rect 220832 4486 220860 200926
rect 221292 180794 221320 200926
rect 222226 200790 222332 200818
rect 222304 200274 222332 200790
rect 222212 200246 222332 200274
rect 222212 197606 222240 200246
rect 222396 200114 222424 200926
rect 222304 200086 222424 200114
rect 222200 197600 222252 197606
rect 222200 197542 222252 197548
rect 220924 180766 221320 180794
rect 220924 6118 220952 180766
rect 222304 13122 222332 200086
rect 222856 180794 222884 200926
rect 223488 198348 223540 198354
rect 223488 198290 223540 198296
rect 222396 180766 222884 180794
rect 222292 13116 222344 13122
rect 222292 13058 222344 13064
rect 222396 9314 222424 180766
rect 222384 9308 222436 9314
rect 222384 9250 222436 9256
rect 220912 6112 220964 6118
rect 220912 6054 220964 6060
rect 221556 5500 221608 5506
rect 221556 5442 221608 5448
rect 220820 4480 220872 4486
rect 220820 4422 220872 4428
rect 221568 480 221596 5442
rect 223500 3398 223528 198290
rect 223684 17270 223712 200926
rect 223960 197402 223988 200926
rect 224512 200114 224540 200926
rect 224144 200086 224540 200114
rect 223948 197396 224000 197402
rect 223948 197338 224000 197344
rect 224144 180794 224172 200086
rect 225064 197810 225092 200926
rect 225052 197804 225104 197810
rect 225052 197746 225104 197752
rect 224224 197600 224276 197606
rect 224224 197542 224276 197548
rect 223868 180766 224172 180794
rect 223672 17264 223724 17270
rect 223672 17206 223724 17212
rect 223868 9382 223896 180766
rect 223856 9376 223908 9382
rect 223856 9318 223908 9324
rect 224236 4214 224264 197542
rect 225432 180794 225460 200926
rect 226366 200790 226472 200818
rect 225064 180766 225460 180794
rect 225064 84930 225092 180766
rect 225052 84924 225104 84930
rect 225052 84866 225104 84872
rect 226444 16046 226472 200790
rect 226536 198490 226564 200926
rect 226524 198484 226576 198490
rect 226524 198426 226576 198432
rect 226996 180794 227024 200926
rect 227732 198558 227760 200926
rect 228008 200114 228036 200926
rect 227824 200086 228036 200114
rect 227720 198552 227772 198558
rect 227720 198494 227772 198500
rect 227628 198416 227680 198422
rect 227628 198358 227680 198364
rect 226536 180766 227024 180794
rect 226432 16040 226484 16046
rect 226432 15982 226484 15988
rect 226536 6050 226564 180766
rect 227640 6914 227668 198358
rect 227824 17474 227852 200086
rect 228560 180794 228588 200926
rect 228008 180766 228588 180794
rect 227812 17468 227864 17474
rect 227812 17410 227864 17416
rect 227548 6886 227668 6914
rect 226524 6044 226576 6050
rect 226524 5986 226576 5992
rect 224224 4208 224276 4214
rect 224224 4150 224276 4156
rect 225144 3936 225196 3942
rect 225144 3878 225196 3884
rect 223948 3800 224000 3806
rect 223948 3742 224000 3748
rect 222752 3392 222804 3398
rect 222752 3334 222804 3340
rect 223488 3392 223540 3398
rect 223488 3334 223540 3340
rect 222764 480 222792 3334
rect 223960 480 223988 3742
rect 225156 480 225184 3878
rect 226340 3664 226392 3670
rect 226340 3606 226392 3612
rect 226352 480 226380 3606
rect 227548 480 227576 6886
rect 228008 5982 228036 180766
rect 229204 13190 229232 200926
rect 229664 198626 229692 200926
rect 230506 200790 230612 200818
rect 229652 198620 229704 198626
rect 229652 198562 229704 198568
rect 229192 13184 229244 13190
rect 229192 13126 229244 13132
rect 227996 5976 228048 5982
rect 227996 5918 228048 5924
rect 230584 5914 230612 200790
rect 230676 7274 230704 200926
rect 231136 180794 231164 200926
rect 231768 198484 231820 198490
rect 231768 198426 231820 198432
rect 230768 180766 231164 180794
rect 230664 7268 230716 7274
rect 230664 7210 230716 7216
rect 230572 5908 230624 5914
rect 230572 5850 230624 5856
rect 230768 4418 230796 180766
rect 230756 4412 230808 4418
rect 230756 4354 230808 4360
rect 228732 4072 228784 4078
rect 228732 4014 228784 4020
rect 228744 480 228772 4014
rect 229836 3732 229888 3738
rect 229836 3674 229888 3680
rect 229848 480 229876 3674
rect 231780 3398 231808 198426
rect 231860 191140 231912 191146
rect 231860 191082 231912 191088
rect 231872 4350 231900 191082
rect 231964 5846 231992 200926
rect 232148 7206 232176 200926
rect 232504 197804 232556 197810
rect 232504 197746 232556 197752
rect 232136 7200 232188 7206
rect 232136 7142 232188 7148
rect 231952 5840 232004 5846
rect 231952 5782 232004 5788
rect 231860 4344 231912 4350
rect 231860 4286 231912 4292
rect 232228 4004 232280 4010
rect 232228 3946 232280 3952
rect 231032 3392 231084 3398
rect 231032 3334 231084 3340
rect 231768 3392 231820 3398
rect 231768 3334 231820 3340
rect 231044 480 231072 3334
rect 232240 480 232268 3946
rect 232516 3874 232544 197746
rect 232792 191146 232820 200926
rect 232780 191140 232832 191146
rect 232780 191082 232832 191088
rect 233252 5778 233280 200926
rect 233712 180794 233740 200926
rect 234646 200790 234752 200818
rect 234724 200114 234752 200790
rect 234632 200086 234752 200114
rect 234528 198552 234580 198558
rect 234528 198494 234580 198500
rect 233344 180766 233740 180794
rect 233344 7138 233372 180766
rect 233332 7132 233384 7138
rect 233332 7074 233384 7080
rect 233240 5772 233292 5778
rect 233240 5714 233292 5720
rect 232504 3868 232556 3874
rect 232504 3810 232556 3816
rect 234540 3398 234568 198494
rect 234632 4282 234660 200086
rect 234816 195242 234844 200926
rect 234724 195214 234844 195242
rect 234724 5710 234752 195214
rect 235276 180794 235304 200926
rect 235908 198620 235960 198626
rect 235908 198562 235960 198568
rect 234816 180766 235304 180794
rect 234816 7070 234844 180766
rect 234804 7064 234856 7070
rect 234804 7006 234856 7012
rect 234712 5704 234764 5710
rect 234712 5646 234764 5652
rect 234620 4276 234672 4282
rect 234620 4218 234672 4224
rect 233424 3392 233476 3398
rect 233424 3334 233476 3340
rect 234528 3392 234580 3398
rect 234528 3334 234580 3340
rect 235816 3392 235868 3398
rect 235816 3334 235868 3340
rect 233436 480 233464 3334
rect 234620 3324 234672 3330
rect 234620 3266 234672 3272
rect 234632 480 234660 3266
rect 235828 480 235856 3334
rect 235920 3330 235948 198562
rect 236012 197674 236040 200926
rect 236288 197742 236316 200926
rect 236276 197736 236328 197742
rect 236276 197678 236328 197684
rect 236000 197668 236052 197674
rect 236000 197610 236052 197616
rect 236748 180794 236776 200926
rect 237380 195288 237432 195294
rect 237380 195230 237432 195236
rect 236288 180766 236776 180794
rect 236288 5642 236316 180766
rect 237392 14686 237420 195230
rect 237484 16114 237512 200926
rect 237944 195294 237972 200926
rect 238786 200790 238892 200818
rect 238668 198688 238720 198694
rect 238668 198630 238720 198636
rect 237932 195288 237984 195294
rect 237932 195230 237984 195236
rect 237472 16108 237524 16114
rect 237472 16050 237524 16056
rect 237380 14680 237432 14686
rect 237380 14622 237432 14628
rect 238024 14544 238076 14550
rect 238024 14486 238076 14492
rect 236276 5636 236328 5642
rect 236276 5578 236328 5584
rect 238036 3942 238064 14486
rect 238024 3936 238076 3942
rect 238024 3878 238076 3884
rect 237012 3868 237064 3874
rect 237012 3810 237064 3816
rect 235908 3324 235960 3330
rect 235908 3266 235960 3272
rect 237024 480 237052 3810
rect 238680 3330 238708 198630
rect 238864 180794 238892 200790
rect 238956 196858 238984 200926
rect 239416 197878 239444 200926
rect 240350 200790 240456 200818
rect 240232 200456 240284 200462
rect 240232 200398 240284 200404
rect 239404 197872 239456 197878
rect 239404 197814 239456 197820
rect 238944 196852 238996 196858
rect 238944 196794 238996 196800
rect 238772 180766 238892 180794
rect 238772 6186 238800 180766
rect 240244 9518 240272 200398
rect 240428 180794 240456 200790
rect 240520 200462 240548 200926
rect 240508 200456 240560 200462
rect 240508 200398 240560 200404
rect 241072 197946 241100 200926
rect 241060 197940 241112 197946
rect 241060 197882 241112 197888
rect 241428 197940 241480 197946
rect 241428 197882 241480 197888
rect 240336 180766 240456 180794
rect 240232 9512 240284 9518
rect 240232 9454 240284 9460
rect 240336 6254 240364 180766
rect 240324 6248 240376 6254
rect 240324 6190 240376 6196
rect 238760 6180 238812 6186
rect 238760 6122 238812 6128
rect 241440 3534 241468 197882
rect 241532 4826 241560 200926
rect 241992 180794 242020 200926
rect 242926 200790 243032 200818
rect 243004 196926 243032 200790
rect 243096 197606 243124 200926
rect 243084 197600 243136 197606
rect 243084 197542 243136 197548
rect 242992 196920 243044 196926
rect 242992 196862 243044 196868
rect 243648 196654 243676 200926
rect 244490 200790 244596 200818
rect 244568 200114 244596 200790
rect 244476 200086 244596 200114
rect 243636 196648 243688 196654
rect 243636 196590 243688 196596
rect 244280 193316 244332 193322
rect 244280 193258 244332 193264
rect 241624 180766 242020 180794
rect 241624 9586 241652 180766
rect 242164 87644 242216 87650
rect 242164 87586 242216 87592
rect 241612 9580 241664 9586
rect 241612 9522 241664 9528
rect 241520 4820 241572 4826
rect 241520 4762 241572 4768
rect 242176 4078 242204 87586
rect 242900 4140 242952 4146
rect 242900 4082 242952 4088
rect 242164 4072 242216 4078
rect 242164 4014 242216 4020
rect 241704 3936 241756 3942
rect 241704 3878 241756 3884
rect 240508 3528 240560 3534
rect 240508 3470 240560 3476
rect 241428 3528 241480 3534
rect 241428 3470 241480 3476
rect 238116 3324 238168 3330
rect 238116 3266 238168 3272
rect 238668 3324 238720 3330
rect 238668 3266 238720 3272
rect 238128 480 238156 3266
rect 239312 3256 239364 3262
rect 239312 3198 239364 3204
rect 239324 480 239352 3198
rect 240520 480 240548 3470
rect 241716 480 241744 3878
rect 242912 480 242940 4082
rect 244096 4072 244148 4078
rect 244096 4014 244148 4020
rect 244108 480 244136 4014
rect 244292 3466 244320 193258
rect 244372 190936 244424 190942
rect 244372 190878 244424 190884
rect 244384 17338 244412 190878
rect 244476 155242 244504 200086
rect 244660 193322 244688 200926
rect 244924 197396 244976 197402
rect 244924 197338 244976 197344
rect 244648 193316 244700 193322
rect 244648 193258 244700 193264
rect 244464 155236 244516 155242
rect 244464 155178 244516 155184
rect 244372 17332 244424 17338
rect 244372 17274 244424 17280
rect 244936 3602 244964 197338
rect 245120 190942 245148 200926
rect 245752 194540 245804 194546
rect 245752 194482 245804 194488
rect 245108 190936 245160 190942
rect 245108 190878 245160 190884
rect 245016 22908 245068 22914
rect 245016 22850 245068 22856
rect 244924 3596 244976 3602
rect 244924 3538 244976 3544
rect 244280 3460 244332 3466
rect 244280 3402 244332 3408
rect 245028 3330 245056 22850
rect 245764 14482 245792 194482
rect 245752 14476 245804 14482
rect 245752 14418 245804 14424
rect 245856 3398 245884 200926
rect 246224 194546 246252 200926
rect 247066 200790 247172 200818
rect 246304 197668 246356 197674
rect 246304 197610 246356 197616
rect 246212 194540 246264 194546
rect 246212 194482 246264 194488
rect 246316 22846 246344 197610
rect 247144 196722 247172 200790
rect 247132 196716 247184 196722
rect 247132 196658 247184 196664
rect 246304 22840 246356 22846
rect 246304 22782 246356 22788
rect 246948 14476 247000 14482
rect 246948 14418 247000 14424
rect 246960 3534 246988 14418
rect 247236 6322 247264 200926
rect 247696 197402 247724 200926
rect 247684 197396 247736 197402
rect 247684 197338 247736 197344
rect 247224 6316 247276 6322
rect 247224 6258 247276 6264
rect 248432 4894 248460 200926
rect 248708 200114 248736 200926
rect 248524 200086 248736 200114
rect 248524 6390 248552 200086
rect 249168 180794 249196 200926
rect 248708 180766 249196 180794
rect 248708 15910 248736 180766
rect 248696 15904 248748 15910
rect 248696 15846 248748 15852
rect 248512 6384 248564 6390
rect 248512 6326 248564 6332
rect 249812 4962 249840 200926
rect 250180 180794 250208 200926
rect 251206 200790 251404 200818
rect 250444 197396 250496 197402
rect 250444 197338 250496 197344
rect 249904 180766 250208 180794
rect 249904 6458 249932 180766
rect 250456 22778 250484 197338
rect 251272 195288 251324 195294
rect 251272 195230 251324 195236
rect 250444 22772 250496 22778
rect 250444 22714 250496 22720
rect 251088 13116 251140 13122
rect 251088 13058 251140 13064
rect 249892 6452 249944 6458
rect 249892 6394 249944 6400
rect 249800 4956 249852 4962
rect 249800 4898 249852 4904
rect 248420 4888 248472 4894
rect 248420 4830 248472 4836
rect 246396 3528 246448 3534
rect 246396 3470 246448 3476
rect 246948 3528 247000 3534
rect 246948 3470 247000 3476
rect 247592 3528 247644 3534
rect 247592 3470 247644 3476
rect 245844 3392 245896 3398
rect 245844 3334 245896 3340
rect 245016 3324 245068 3330
rect 245016 3266 245068 3272
rect 245200 3324 245252 3330
rect 245200 3266 245252 3272
rect 245212 480 245240 3266
rect 246408 480 246436 3470
rect 247604 480 247632 3470
rect 251100 3466 251128 13058
rect 251284 6526 251312 195230
rect 251376 84998 251404 200790
rect 251364 84992 251416 84998
rect 251364 84934 251416 84940
rect 251272 6520 251324 6526
rect 251272 6462 251324 6468
rect 251468 5030 251496 200926
rect 251824 197736 251876 197742
rect 251824 197678 251876 197684
rect 251456 5024 251508 5030
rect 251456 4966 251508 4972
rect 251180 3596 251232 3602
rect 251180 3538 251232 3544
rect 249984 3460 250036 3466
rect 249984 3402 250036 3408
rect 251088 3460 251140 3466
rect 251088 3402 251140 3408
rect 248788 3120 248840 3126
rect 248788 3062 248840 3068
rect 248800 480 248828 3062
rect 249996 480 250024 3402
rect 251192 480 251220 3538
rect 251836 3330 251864 197678
rect 251928 195294 251956 200926
rect 252678 200790 252784 200818
rect 252560 200456 252612 200462
rect 252560 200398 252612 200404
rect 251916 195288 251968 195294
rect 251916 195230 251968 195236
rect 252572 4758 252600 200398
rect 252756 86290 252784 200790
rect 252848 200462 252876 200926
rect 252836 200456 252888 200462
rect 252836 200398 252888 200404
rect 253308 180794 253336 200926
rect 253848 197872 253900 197878
rect 253848 197814 253900 197820
rect 252848 180766 253336 180794
rect 252744 86284 252796 86290
rect 252744 86226 252796 86232
rect 252848 6594 252876 180766
rect 252836 6588 252888 6594
rect 252836 6530 252888 6536
rect 252560 4752 252612 4758
rect 252560 4694 252612 4700
rect 251824 3324 251876 3330
rect 251824 3266 251876 3272
rect 252376 3052 252428 3058
rect 252376 2994 252428 3000
rect 252388 480 252416 2994
rect 253492 598 253704 626
rect 253492 480 253520 598
rect 253676 490 253704 598
rect 253860 490 253888 197814
rect 253952 197402 253980 200926
rect 253940 197396 253992 197402
rect 253940 197338 253992 197344
rect 254032 195288 254084 195294
rect 254032 195230 254084 195236
rect 254044 6662 254072 195230
rect 254320 180794 254348 200926
rect 254872 195294 254900 200926
rect 255424 198014 255452 200926
rect 255412 198008 255464 198014
rect 255412 197950 255464 197956
rect 254860 195288 254912 195294
rect 254860 195230 254912 195236
rect 255884 180794 255912 200926
rect 256818 200790 256924 200818
rect 256896 200114 256924 200790
rect 256804 200086 256924 200114
rect 255964 198008 256016 198014
rect 255964 197950 256016 197956
rect 254136 180766 254348 180794
rect 255424 180766 255912 180794
rect 254032 6656 254084 6662
rect 254032 6598 254084 6604
rect 254136 4690 254164 180766
rect 255424 5234 255452 180766
rect 255412 5228 255464 5234
rect 255412 5170 255464 5176
rect 254124 4684 254176 4690
rect 254124 4626 254176 4632
rect 254676 3392 254728 3398
rect 254676 3334 254728 3340
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9926 -960 10038 480
rect 11122 -960 11234 480
rect 12318 -960 12430 480
rect 13514 -960 13626 480
rect 14710 -960 14822 480
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 18206 -960 18318 480
rect 19402 -960 19514 480
rect 20598 -960 20710 480
rect 21794 -960 21906 480
rect 22990 -960 23102 480
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26486 -960 26598 480
rect 27682 -960 27794 480
rect 28878 -960 28990 480
rect 30074 -960 30186 480
rect 31270 -960 31382 480
rect 32374 -960 32486 480
rect 33570 -960 33682 480
rect 34766 -960 34878 480
rect 35962 -960 36074 480
rect 37158 -960 37270 480
rect 38354 -960 38466 480
rect 39550 -960 39662 480
rect 40654 -960 40766 480
rect 41850 -960 41962 480
rect 43046 -960 43158 480
rect 44242 -960 44354 480
rect 45438 -960 45550 480
rect 46634 -960 46746 480
rect 47830 -960 47942 480
rect 48934 -960 49046 480
rect 50130 -960 50242 480
rect 51326 -960 51438 480
rect 52522 -960 52634 480
rect 53718 -960 53830 480
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 57214 -960 57326 480
rect 58410 -960 58522 480
rect 59606 -960 59718 480
rect 60802 -960 60914 480
rect 61998 -960 62110 480
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65494 -960 65606 480
rect 66690 -960 66802 480
rect 67886 -960 67998 480
rect 69082 -960 69194 480
rect 70278 -960 70390 480
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73774 -960 73886 480
rect 74970 -960 75082 480
rect 76166 -960 76278 480
rect 77362 -960 77474 480
rect 78558 -960 78670 480
rect 79662 -960 79774 480
rect 80858 -960 80970 480
rect 82054 -960 82166 480
rect 83250 -960 83362 480
rect 84446 -960 84558 480
rect 85642 -960 85754 480
rect 86838 -960 86950 480
rect 87942 -960 88054 480
rect 89138 -960 89250 480
rect 90334 -960 90446 480
rect 91530 -960 91642 480
rect 92726 -960 92838 480
rect 93922 -960 94034 480
rect 95118 -960 95230 480
rect 96222 -960 96334 480
rect 97418 -960 97530 480
rect 98614 -960 98726 480
rect 99810 -960 99922 480
rect 101006 -960 101118 480
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104502 -960 104614 480
rect 105698 -960 105810 480
rect 106894 -960 107006 480
rect 108090 -960 108202 480
rect 109286 -960 109398 480
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112782 -960 112894 480
rect 113978 -960 114090 480
rect 115174 -960 115286 480
rect 116370 -960 116482 480
rect 117566 -960 117678 480
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 121062 -960 121174 480
rect 122258 -960 122370 480
rect 123454 -960 123566 480
rect 124650 -960 124762 480
rect 125846 -960 125958 480
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 129342 -960 129454 480
rect 130538 -960 130650 480
rect 131734 -960 131846 480
rect 132930 -960 133042 480
rect 134126 -960 134238 480
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137622 -960 137734 480
rect 138818 -960 138930 480
rect 140014 -960 140126 480
rect 141210 -960 141322 480
rect 142406 -960 142518 480
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145902 -960 146014 480
rect 147098 -960 147210 480
rect 148294 -960 148406 480
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 154182 -960 154294 480
rect 155378 -960 155490 480
rect 156574 -960 156686 480
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162462 -960 162574 480
rect 163658 -960 163770 480
rect 164854 -960 164966 480
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170742 -960 170854 480
rect 171938 -960 172050 480
rect 173134 -960 173246 480
rect 174238 -960 174350 480
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 179022 -960 179134 480
rect 180218 -960 180330 480
rect 181414 -960 181526 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 187302 -960 187414 480
rect 188498 -960 188610 480
rect 189694 -960 189806 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 199078 -960 199190 480
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207358 -960 207470 480
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 212142 -960 212254 480
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215638 -960 215750 480
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220422 -960 220534 480
rect 221526 -960 221638 480
rect 222722 -960 222834 480
rect 223918 -960 224030 480
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228702 -960 228814 480
rect 229806 -960 229918 480
rect 231002 -960 231114 480
rect 232198 -960 232310 480
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236982 -960 237094 480
rect 238086 -960 238198 480
rect 239282 -960 239394 480
rect 240478 -960 240590 480
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 246366 -960 246478 480
rect 247562 -960 247674 480
rect 248758 -960 248870 480
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 253676 462 253888 490
rect 254688 480 254716 3334
rect 255872 3324 255924 3330
rect 255872 3266 255924 3272
rect 255884 480 255912 3266
rect 255976 3058 256004 197950
rect 256056 197532 256108 197538
rect 256056 197474 256108 197480
rect 256068 3806 256096 197474
rect 256804 177342 256832 200086
rect 257080 198082 257108 200926
rect 257068 198076 257120 198082
rect 257068 198018 257120 198024
rect 257448 180794 257476 200926
rect 256896 180766 257476 180794
rect 256792 177336 256844 177342
rect 256792 177278 256844 177284
rect 256896 5302 256924 180766
rect 258184 171834 258212 200926
rect 258552 198150 258580 200926
rect 258540 198144 258592 198150
rect 258540 198086 258592 198092
rect 259012 180794 259040 200926
rect 259368 198076 259420 198082
rect 259368 198018 259420 198024
rect 258276 180766 259040 180794
rect 258172 171828 258224 171834
rect 258172 171770 258224 171776
rect 258276 5370 258304 180766
rect 258724 176724 258776 176730
rect 258724 176666 258776 176672
rect 258264 5364 258316 5370
rect 258264 5306 258316 5312
rect 256884 5296 256936 5302
rect 256884 5238 256936 5244
rect 256056 3800 256108 3806
rect 256056 3742 256108 3748
rect 258736 3670 258764 176666
rect 258264 3664 258316 3670
rect 258184 3612 258264 3618
rect 258184 3606 258316 3612
rect 258724 3664 258776 3670
rect 258724 3606 258776 3612
rect 258184 3590 258304 3606
rect 258184 3466 258212 3590
rect 259380 3466 259408 198018
rect 259656 197674 259684 200926
rect 260208 198218 260236 200926
rect 260958 200790 261064 200818
rect 260196 198212 260248 198218
rect 260196 198154 260248 198160
rect 260656 198144 260708 198150
rect 260656 198086 260708 198092
rect 259644 197668 259696 197674
rect 259644 197610 259696 197616
rect 260104 197532 260156 197538
rect 260104 197474 260156 197480
rect 258172 3460 258224 3466
rect 258172 3402 258224 3408
rect 258264 3460 258316 3466
rect 258264 3402 258316 3408
rect 259368 3460 259420 3466
rect 259368 3402 259420 3408
rect 259460 3460 259512 3466
rect 259460 3402 259512 3408
rect 257068 3188 257120 3194
rect 257068 3130 257120 3136
rect 255964 3052 256016 3058
rect 255964 2994 256016 3000
rect 257080 480 257108 3130
rect 258276 480 258304 3402
rect 259472 480 259500 3402
rect 260116 3262 260144 197474
rect 260668 16574 260696 198086
rect 260748 197668 260800 197674
rect 260748 197610 260800 197616
rect 260576 16546 260696 16574
rect 260576 3466 260604 16546
rect 260760 6914 260788 197610
rect 260668 6886 260788 6914
rect 260564 3460 260616 3466
rect 260564 3402 260616 3408
rect 260104 3256 260156 3262
rect 260104 3198 260156 3204
rect 260668 480 260696 6886
rect 261036 5438 261064 200790
rect 261128 197810 261156 200926
rect 261680 198286 261708 200926
rect 261668 198280 261720 198286
rect 261668 198222 261720 198228
rect 261116 197804 261168 197810
rect 261116 197746 261168 197752
rect 262416 5506 262444 200926
rect 262784 198354 262812 200926
rect 262772 198348 262824 198354
rect 262772 198290 262824 198296
rect 262956 198212 263008 198218
rect 262956 198154 263008 198160
rect 262864 197396 262916 197402
rect 262864 197338 262916 197344
rect 262404 5500 262456 5506
rect 262404 5442 262456 5448
rect 261024 5432 261076 5438
rect 261024 5374 261076 5380
rect 262876 3738 262904 197338
rect 262864 3732 262916 3738
rect 262864 3674 262916 3680
rect 262968 3466 262996 198154
rect 263152 197606 263180 200926
rect 263140 197600 263192 197606
rect 263140 197542 263192 197548
rect 263704 14550 263732 200926
rect 264244 197464 264296 197470
rect 264244 197406 264296 197412
rect 263692 14544 263744 14550
rect 263692 14486 263744 14492
rect 264256 3874 264284 197406
rect 264348 197402 264376 200926
rect 264992 198422 265020 200926
rect 264980 198416 265032 198422
rect 264980 198358 265032 198364
rect 264888 198280 264940 198286
rect 264888 198222 264940 198228
rect 264336 197396 264388 197402
rect 264336 197338 264388 197344
rect 264244 3868 264296 3874
rect 264244 3810 264296 3816
rect 263048 3800 263100 3806
rect 263048 3742 263100 3748
rect 261760 3460 261812 3466
rect 261760 3402 261812 3408
rect 262956 3460 263008 3466
rect 262956 3402 263008 3408
rect 261772 480 261800 3402
rect 263060 1306 263088 3742
rect 264900 3466 264928 198222
rect 265176 87650 265204 200926
rect 265728 197470 265756 200926
rect 266372 198490 266400 200926
rect 266360 198484 266412 198490
rect 266360 198426 266412 198432
rect 265716 197464 265768 197470
rect 265716 197406 265768 197412
rect 266740 180794 266768 200926
rect 267384 198558 267412 200926
rect 267936 198626 267964 200926
rect 267924 198620 267976 198626
rect 267924 198562 267976 198568
rect 267372 198552 267424 198558
rect 267372 198494 267424 198500
rect 267648 198416 267700 198422
rect 267648 198358 267700 198364
rect 267096 197600 267148 197606
rect 267096 197542 267148 197548
rect 267004 197396 267056 197402
rect 267004 197338 267056 197344
rect 266556 180766 266768 180794
rect 266556 176730 266584 180766
rect 266544 176724 266596 176730
rect 266544 176666 266596 176672
rect 265164 87644 265216 87650
rect 265164 87586 265216 87592
rect 267016 4078 267044 197338
rect 267108 4146 267136 197542
rect 267096 4140 267148 4146
rect 267096 4082 267148 4088
rect 267004 4072 267056 4078
rect 267004 4014 267056 4020
rect 265348 3664 265400 3670
rect 265348 3606 265400 3612
rect 264152 3460 264204 3466
rect 264152 3402 264204 3408
rect 264888 3460 264940 3466
rect 264888 3402 264940 3408
rect 262968 1278 263088 1306
rect 262968 480 262996 1278
rect 264164 480 264192 3402
rect 265360 480 265388 3606
rect 267660 3466 267688 198358
rect 268304 180794 268332 200926
rect 269028 198552 269080 198558
rect 269028 198494 269080 198500
rect 268936 198348 268988 198354
rect 268936 198290 268988 198296
rect 268384 197804 268436 197810
rect 268384 197746 268436 197752
rect 267844 180766 268332 180794
rect 267844 22914 267872 180766
rect 267832 22908 267884 22914
rect 267832 22850 267884 22856
rect 266544 3460 266596 3466
rect 266544 3402 266596 3408
rect 267648 3460 267700 3466
rect 267648 3402 267700 3408
rect 266556 480 266584 3402
rect 268396 3194 268424 197746
rect 268948 6914 268976 198290
rect 268856 6886 268976 6914
rect 268384 3188 268436 3194
rect 268384 3130 268436 3136
rect 267740 2916 267792 2922
rect 267740 2858 267792 2864
rect 267752 480 267780 2858
rect 268856 480 268884 6886
rect 269040 2922 269068 198494
rect 269132 197402 269160 200926
rect 269408 198694 269436 200926
rect 269396 198688 269448 198694
rect 269396 198630 269448 198636
rect 269960 197538 269988 200926
rect 270408 198484 270460 198490
rect 270408 198426 270460 198432
rect 269948 197532 270000 197538
rect 269948 197474 270000 197480
rect 269764 197464 269816 197470
rect 269764 197406 269816 197412
rect 269120 197396 269172 197402
rect 269120 197338 269172 197344
rect 269776 4010 269804 197406
rect 269856 197396 269908 197402
rect 269856 197338 269908 197344
rect 269764 4004 269816 4010
rect 269764 3946 269816 3952
rect 269868 3942 269896 197338
rect 269856 3936 269908 3942
rect 269856 3878 269908 3884
rect 269028 2916 269080 2922
rect 269028 2858 269080 2864
rect 270052 598 270264 626
rect 270052 480 270080 598
rect 270236 490 270264 598
rect 270420 490 270448 198426
rect 270604 197946 270632 200926
rect 270592 197940 270644 197946
rect 270592 197882 270644 197888
rect 270880 197402 270908 200926
rect 271432 197606 271460 200926
rect 271788 198620 271840 198626
rect 271788 198562 271840 198568
rect 271420 197600 271472 197606
rect 271420 197542 271472 197548
rect 270868 197396 270920 197402
rect 270868 197338 270920 197344
rect 271144 197396 271196 197402
rect 271144 197338 271196 197344
rect 271156 3534 271184 197338
rect 271800 3534 271828 198562
rect 271984 197470 272012 200926
rect 272536 197742 272564 200926
rect 273378 200790 273484 200818
rect 273456 200114 273484 200790
rect 273364 200086 273484 200114
rect 272524 197736 272576 197742
rect 272524 197678 272576 197684
rect 271972 197464 272024 197470
rect 271972 197406 272024 197412
rect 273364 14482 273392 200086
rect 273640 197402 273668 200926
rect 274008 200114 274036 200926
rect 273824 200086 274036 200114
rect 273628 197396 273680 197402
rect 273628 197338 273680 197344
rect 273824 180794 273852 200086
rect 273904 197396 273956 197402
rect 273904 197338 273956 197344
rect 273456 180766 273852 180794
rect 273352 14476 273404 14482
rect 273352 14418 273404 14424
rect 271144 3528 271196 3534
rect 271144 3470 271196 3476
rect 271236 3528 271288 3534
rect 271236 3470 271288 3476
rect 271788 3528 271840 3534
rect 271788 3470 271840 3476
rect 254646 -960 254758 480
rect 255842 -960 255954 480
rect 257038 -960 257150 480
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262926 -960 263038 480
rect 264122 -960 264234 480
rect 265318 -960 265430 480
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268814 -960 268926 480
rect 270010 -960 270122 480
rect 270236 462 270448 490
rect 271248 480 271276 3470
rect 272432 3392 272484 3398
rect 272432 3334 272484 3340
rect 272444 480 272472 3334
rect 273456 3126 273484 180766
rect 273916 3602 273944 197338
rect 274836 13122 274864 200926
rect 275112 197402 275140 200926
rect 275664 198014 275692 200926
rect 275652 198008 275704 198014
rect 275652 197950 275704 197956
rect 276216 197878 276244 200926
rect 276204 197872 276256 197878
rect 276204 197814 276256 197820
rect 275100 197396 275152 197402
rect 275100 197338 275152 197344
rect 276584 180794 276612 200926
rect 277518 200790 277624 200818
rect 277308 198688 277360 198694
rect 277308 198630 277360 198636
rect 276664 198008 276716 198014
rect 276664 197950 276716 197956
rect 276216 180766 276612 180794
rect 274824 13116 274876 13122
rect 274824 13058 274876 13064
rect 273904 3596 273956 3602
rect 273904 3538 273956 3544
rect 276020 3596 276072 3602
rect 276020 3538 276072 3544
rect 274824 3528 274876 3534
rect 274824 3470 274876 3476
rect 273628 3460 273680 3466
rect 273628 3402 273680 3408
rect 273444 3120 273496 3126
rect 273444 3062 273496 3068
rect 273640 480 273668 3402
rect 274836 480 274864 3470
rect 276032 480 276060 3538
rect 276216 3330 276244 180766
rect 276676 3534 276704 197950
rect 277320 3602 277348 198630
rect 277308 3596 277360 3602
rect 277308 3538 277360 3544
rect 276664 3528 276716 3534
rect 276664 3470 276716 3476
rect 277124 3528 277176 3534
rect 277124 3470 277176 3476
rect 276204 3324 276256 3330
rect 276204 3266 276256 3272
rect 277136 480 277164 3470
rect 277596 3262 277624 200790
rect 277688 197810 277716 200926
rect 278240 198082 278268 200926
rect 278792 198150 278820 200926
rect 278780 198144 278832 198150
rect 278780 198086 278832 198092
rect 278228 198076 278280 198082
rect 278228 198018 278280 198024
rect 278688 198076 278740 198082
rect 278688 198018 278740 198024
rect 277676 197804 277728 197810
rect 277676 197746 277728 197752
rect 277584 3256 277636 3262
rect 277584 3198 277636 3204
rect 278332 598 278544 626
rect 278332 480 278360 598
rect 278516 490 278544 598
rect 278700 490 278728 198018
rect 279160 197674 279188 200926
rect 279712 198218 279740 200926
rect 279700 198212 279752 198218
rect 279700 198154 279752 198160
rect 279148 197668 279200 197674
rect 279148 197610 279200 197616
rect 280356 3806 280384 200926
rect 280816 198286 280844 200926
rect 280804 198280 280856 198286
rect 280804 198222 280856 198228
rect 281552 197402 281580 200926
rect 281736 198422 281764 200926
rect 282288 198558 282316 200926
rect 282276 198552 282328 198558
rect 282276 198494 282328 198500
rect 281724 198416 281776 198422
rect 281724 198358 281776 198364
rect 282932 198354 282960 200926
rect 283392 198490 283420 200926
rect 283944 198626 283972 200926
rect 283932 198620 283984 198626
rect 283932 198562 283984 198568
rect 283380 198484 283432 198490
rect 283380 198426 283432 198432
rect 282920 198348 282972 198354
rect 282920 198290 282972 198296
rect 282184 197464 282236 197470
rect 282184 197406 282236 197412
rect 280804 197396 280856 197402
rect 280804 197338 280856 197344
rect 281540 197396 281592 197402
rect 281540 197338 281592 197344
rect 280344 3800 280396 3806
rect 280344 3742 280396 3748
rect 280816 3670 280844 197338
rect 281908 4140 281960 4146
rect 281908 4082 281960 4088
rect 280804 3664 280856 3670
rect 280804 3606 280856 3612
rect 279516 3596 279568 3602
rect 279516 3538 279568 3544
rect 271206 -960 271318 480
rect 272402 -960 272514 480
rect 273598 -960 273710 480
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 277094 -960 277206 480
rect 278290 -960 278402 480
rect 278516 462 278728 490
rect 279528 480 279556 3538
rect 280712 3324 280764 3330
rect 280712 3266 280764 3272
rect 280724 480 280752 3266
rect 281920 480 281948 4082
rect 282196 3466 282224 197406
rect 284312 197402 284340 200926
rect 284864 197470 284892 200926
rect 285588 198280 285640 198286
rect 285588 198222 285640 198228
rect 285496 198144 285548 198150
rect 285496 198086 285548 198092
rect 284852 197464 284904 197470
rect 284852 197406 284904 197412
rect 284944 197464 284996 197470
rect 284944 197406 284996 197412
rect 282276 197396 282328 197402
rect 282276 197338 282328 197344
rect 284300 197396 284352 197402
rect 284300 197338 284352 197344
rect 282184 3460 282236 3466
rect 282184 3402 282236 3408
rect 282288 3398 282316 197338
rect 284300 3664 284352 3670
rect 284300 3606 284352 3612
rect 282276 3392 282328 3398
rect 282276 3334 282328 3340
rect 283104 3120 283156 3126
rect 283104 3062 283156 3068
rect 283116 480 283144 3062
rect 284312 480 284340 3606
rect 284956 3534 284984 197406
rect 285508 3670 285536 198086
rect 285496 3664 285548 3670
rect 285496 3606 285548 3612
rect 284944 3528 284996 3534
rect 285600 3516 285628 198222
rect 285692 198014 285720 200926
rect 285968 198694 285996 200926
rect 285956 198688 286008 198694
rect 285956 198630 286008 198636
rect 285680 198008 285732 198014
rect 285680 197950 285732 197956
rect 286520 197470 286548 200926
rect 287072 198082 287100 200926
rect 287060 198076 287112 198082
rect 287060 198018 287112 198024
rect 286968 198008 287020 198014
rect 286968 197950 287020 197956
rect 286508 197464 286560 197470
rect 286508 197406 286560 197412
rect 286324 197396 286376 197402
rect 286324 197338 286376 197344
rect 286336 3602 286364 197338
rect 286324 3596 286376 3602
rect 286324 3538 286376 3544
rect 284944 3470 284996 3476
rect 285416 3488 285628 3516
rect 285416 480 285444 3488
rect 286612 598 286824 626
rect 286612 480 286640 598
rect 286796 490 286824 598
rect 286980 490 287008 197950
rect 287440 197402 287468 200926
rect 287900 200114 287928 200926
rect 287624 200086 287928 200114
rect 287428 197396 287480 197402
rect 287428 197338 287480 197344
rect 287624 180794 287652 200086
rect 287704 197396 287756 197402
rect 287704 197338 287756 197344
rect 287348 180766 287652 180794
rect 287348 3330 287376 180766
rect 287336 3324 287388 3330
rect 287336 3266 287388 3272
rect 287716 3126 287744 197338
rect 288544 4146 288572 200926
rect 289096 197402 289124 200926
rect 289832 198150 289860 200926
rect 290108 198286 290136 200926
rect 290096 198280 290148 198286
rect 290096 198222 290148 198228
rect 289820 198144 289872 198150
rect 289820 198086 289872 198092
rect 290568 198014 290596 200926
rect 290556 198008 290608 198014
rect 290556 197950 290608 197956
rect 289084 197396 289136 197402
rect 289084 197338 289136 197344
rect 289728 197396 289780 197402
rect 289728 197338 289780 197344
rect 288532 4140 288584 4146
rect 288532 4082 288584 4088
rect 289740 3534 289768 197338
rect 288992 3528 289044 3534
rect 288992 3470 289044 3476
rect 289728 3528 289780 3534
rect 289728 3470 289780 3476
rect 287796 3188 287848 3194
rect 287796 3130 287848 3136
rect 287704 3120 287756 3126
rect 287704 3062 287756 3068
rect 279486 -960 279598 480
rect 280682 -960 280794 480
rect 281878 -960 281990 480
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 285374 -960 285486 480
rect 286570 -960 286682 480
rect 286796 462 287008 490
rect 287808 480 287836 3130
rect 289004 480 289032 3470
rect 291304 3194 291332 200926
rect 291672 197402 291700 200926
rect 291660 197396 291712 197402
rect 291660 197338 291712 197344
rect 292132 180794 292160 200926
rect 292592 197418 292620 200926
rect 291488 180766 292160 180794
rect 292500 197390 292620 197418
rect 291384 3528 291436 3534
rect 291384 3470 291436 3476
rect 291292 3188 291344 3194
rect 291292 3130 291344 3136
rect 290188 2984 290240 2990
rect 290188 2926 290240 2932
rect 290200 480 290228 2926
rect 291396 480 291424 3470
rect 291488 2990 291516 180766
rect 292500 3534 292528 197390
rect 293052 180794 293080 200926
rect 293986 200790 294092 200818
rect 294064 200114 294092 200790
rect 292776 180766 293080 180794
rect 293972 200086 294092 200114
rect 292776 6914 292804 180766
rect 292592 6886 292804 6914
rect 292488 3528 292540 3534
rect 292488 3470 292540 3476
rect 291476 2984 291528 2990
rect 291476 2926 291528 2932
rect 292592 480 292620 6886
rect 293972 2802 294000 200086
rect 294248 180794 294276 200926
rect 295090 200790 295288 200818
rect 295550 200790 295840 200818
rect 296102 200790 296392 200818
rect 296562 200790 296668 200818
rect 297114 200790 297496 200818
rect 297666 200790 298048 200818
rect 298126 200790 298416 200818
rect 298678 200790 298968 200818
rect 299230 200790 299336 200818
rect 299690 200790 300072 200818
rect 300242 200790 300624 200818
rect 300702 200790 300808 200818
rect 301254 200790 301544 200818
rect 301806 200790 302096 200818
rect 302266 200790 302648 200818
rect 302818 200790 303200 200818
rect 303278 200790 303568 200818
rect 303830 200790 304120 200818
rect 304382 200790 304672 200818
rect 304842 200790 304948 200818
rect 305394 200790 305776 200818
rect 305946 200790 306328 200818
rect 306406 200790 306696 200818
rect 306958 200790 307248 200818
rect 307418 200790 307616 200818
rect 307970 200790 308352 200818
rect 308522 200790 308904 200818
rect 308982 200790 309088 200818
rect 309534 200790 309824 200818
rect 309994 200790 310376 200818
rect 310546 200790 310928 200818
rect 311098 200790 311480 200818
rect 311558 200790 311848 200818
rect 312110 200790 312400 200818
rect 312570 200790 312952 200818
rect 313122 200790 313228 200818
rect 313674 200790 314056 200818
rect 314134 200790 314516 200818
rect 314686 200790 314976 200818
rect 315238 200790 315528 200818
rect 315698 200790 315988 200818
rect 316250 200790 316632 200818
rect 316710 200790 317184 200818
rect 317262 200790 317368 200818
rect 317814 200790 318012 200818
rect 318274 200790 318564 200818
rect 318826 200790 319208 200818
rect 319286 200790 319576 200818
rect 319838 200790 320128 200818
rect 320390 200790 320680 200818
rect 320850 200790 321140 200818
rect 295260 197418 295288 200790
rect 295812 198014 295840 200790
rect 295800 198008 295852 198014
rect 295800 197950 295852 197956
rect 296364 197538 296392 200790
rect 296640 200114 296668 200790
rect 296548 200086 296668 200114
rect 296352 197532 296404 197538
rect 296352 197474 296404 197480
rect 295260 197390 295380 197418
rect 295352 190454 295380 197390
rect 295352 190426 295564 190454
rect 294064 180766 294276 180794
rect 294064 3534 294092 180766
rect 295536 16574 295564 190426
rect 295536 16546 295656 16574
rect 294052 3528 294104 3534
rect 294052 3470 294104 3476
rect 294880 3528 294932 3534
rect 294880 3470 294932 3476
rect 293696 2774 294000 2802
rect 293696 480 293724 2774
rect 294892 480 294920 3470
rect 295628 490 295656 16546
rect 296548 3466 296576 200086
rect 296628 198008 296680 198014
rect 296628 197950 296680 197956
rect 296640 4146 296668 197950
rect 297468 197402 297496 200790
rect 298020 197878 298048 200790
rect 298388 198558 298416 200790
rect 298376 198552 298428 198558
rect 298376 198494 298428 198500
rect 298008 197872 298060 197878
rect 298008 197814 298060 197820
rect 298744 197872 298796 197878
rect 298744 197814 298796 197820
rect 298100 197532 298152 197538
rect 298100 197474 298152 197480
rect 297456 197396 297508 197402
rect 297456 197338 297508 197344
rect 296628 4140 296680 4146
rect 296628 4082 296680 4088
rect 297272 4140 297324 4146
rect 297272 4082 297324 4088
rect 296536 3460 296588 3466
rect 296536 3402 296588 3408
rect 295904 598 296116 626
rect 295904 490 295932 598
rect 287766 -960 287878 480
rect 288962 -960 289074 480
rect 290158 -960 290270 480
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293654 -960 293766 480
rect 294850 -960 294962 480
rect 295628 462 295932 490
rect 296088 480 296116 598
rect 297284 480 297312 4082
rect 298112 490 298140 197474
rect 298756 3194 298784 197814
rect 298940 197402 298968 200790
rect 299308 198422 299336 200790
rect 299296 198416 299348 198422
rect 299296 198358 299348 198364
rect 300044 197470 300072 200790
rect 300596 200114 300624 200790
rect 300596 200086 300716 200114
rect 300032 197464 300084 197470
rect 300032 197406 300084 197412
rect 298836 197396 298888 197402
rect 298836 197338 298888 197344
rect 298928 197396 298980 197402
rect 298928 197338 298980 197344
rect 300124 197396 300176 197402
rect 300124 197338 300176 197344
rect 298744 3188 298796 3194
rect 298744 3130 298796 3136
rect 298848 3058 298876 197338
rect 300136 3534 300164 197338
rect 300688 3874 300716 200086
rect 300780 197606 300808 200790
rect 300768 197600 300820 197606
rect 300768 197542 300820 197548
rect 301516 197470 301544 200790
rect 302068 197538 302096 200790
rect 302516 198552 302568 198558
rect 302516 198494 302568 198500
rect 302056 197532 302108 197538
rect 302056 197474 302108 197480
rect 300768 197464 300820 197470
rect 300768 197406 300820 197412
rect 301504 197464 301556 197470
rect 301504 197406 301556 197412
rect 300780 3942 300808 197406
rect 302528 16574 302556 198494
rect 302620 198082 302648 200790
rect 303172 200114 303200 200790
rect 303172 200086 303476 200114
rect 302608 198076 302660 198082
rect 302608 198018 302660 198024
rect 302528 16546 303200 16574
rect 300768 3936 300820 3942
rect 300768 3878 300820 3884
rect 300676 3868 300728 3874
rect 300676 3810 300728 3816
rect 300124 3528 300176 3534
rect 300124 3470 300176 3476
rect 299664 3460 299716 3466
rect 299664 3402 299716 3408
rect 298836 3052 298888 3058
rect 298836 2994 298888 3000
rect 298296 598 298508 626
rect 298296 490 298324 598
rect 296046 -960 296158 480
rect 297242 -960 297354 480
rect 298112 462 298324 490
rect 298480 480 298508 598
rect 299676 480 299704 3402
rect 301964 3188 302016 3194
rect 301964 3130 302016 3136
rect 300768 3052 300820 3058
rect 300768 2994 300820 3000
rect 300780 480 300808 2994
rect 301976 480 302004 3130
rect 303172 480 303200 16546
rect 303448 4146 303476 200086
rect 303436 4140 303488 4146
rect 303436 4082 303488 4088
rect 303540 3602 303568 200790
rect 304092 198218 304120 200790
rect 304644 200114 304672 200790
rect 304644 200086 304856 200114
rect 304080 198212 304132 198218
rect 304080 198154 304132 198160
rect 304264 197532 304316 197538
rect 304264 197474 304316 197480
rect 303528 3596 303580 3602
rect 303528 3538 303580 3544
rect 304276 3398 304304 197474
rect 304356 3528 304408 3534
rect 304356 3470 304408 3476
rect 304264 3392 304316 3398
rect 304264 3334 304316 3340
rect 304368 480 304396 3470
rect 304828 3466 304856 200086
rect 304920 3806 304948 200790
rect 305184 198416 305236 198422
rect 305184 198358 305236 198364
rect 305196 16574 305224 198358
rect 305644 197600 305696 197606
rect 305644 197542 305696 197548
rect 305196 16546 305592 16574
rect 304908 3800 304960 3806
rect 304908 3742 304960 3748
rect 304816 3460 304868 3466
rect 304816 3402 304868 3408
rect 305564 480 305592 16546
rect 305656 3670 305684 197542
rect 305748 197402 305776 200790
rect 305736 197396 305788 197402
rect 305736 197338 305788 197344
rect 306196 197396 306248 197402
rect 306196 197338 306248 197344
rect 306208 4078 306236 197338
rect 306196 4072 306248 4078
rect 306196 4014 306248 4020
rect 306300 4010 306328 200790
rect 306668 197742 306696 200790
rect 307220 198014 307248 200790
rect 307208 198008 307260 198014
rect 307208 197950 307260 197956
rect 306656 197736 306708 197742
rect 306656 197678 306708 197684
rect 307024 197464 307076 197470
rect 307024 197406 307076 197412
rect 306288 4004 306340 4010
rect 306288 3946 306340 3952
rect 306748 3936 306800 3942
rect 306748 3878 306800 3884
rect 305644 3664 305696 3670
rect 305644 3606 305696 3612
rect 306760 480 306788 3878
rect 307036 3194 307064 197406
rect 307588 5302 307616 200790
rect 307668 197736 307720 197742
rect 307668 197678 307720 197684
rect 307576 5296 307628 5302
rect 307576 5238 307628 5244
rect 307680 3602 307708 197678
rect 308324 197402 308352 200790
rect 308312 197396 308364 197402
rect 308312 197338 308364 197344
rect 308876 190454 308904 200790
rect 309060 197606 309088 200790
rect 309796 198150 309824 200790
rect 309784 198144 309836 198150
rect 309784 198086 309836 198092
rect 310348 197946 310376 200790
rect 310428 198144 310480 198150
rect 310428 198086 310480 198092
rect 310336 197940 310388 197946
rect 310336 197882 310388 197888
rect 309048 197600 309100 197606
rect 309048 197542 309100 197548
rect 309876 197600 309928 197606
rect 309876 197542 309928 197548
rect 309784 197396 309836 197402
rect 309784 197338 309836 197344
rect 308876 190426 309088 190454
rect 309060 6914 309088 190426
rect 308968 6886 309088 6914
rect 307944 3868 307996 3874
rect 307944 3810 307996 3816
rect 307668 3596 307720 3602
rect 307668 3538 307720 3544
rect 307024 3188 307076 3194
rect 307024 3130 307076 3136
rect 307956 480 307984 3810
rect 308968 3738 308996 6886
rect 309796 3874 309824 197338
rect 309888 5234 309916 197542
rect 309876 5228 309928 5234
rect 309876 5170 309928 5176
rect 309784 3868 309836 3874
rect 309784 3810 309836 3816
rect 308956 3732 309008 3738
rect 308956 3674 309008 3680
rect 309048 3664 309100 3670
rect 309048 3606 309100 3612
rect 309060 480 309088 3606
rect 310440 3330 310468 198086
rect 310900 197742 310928 200790
rect 311452 200114 311480 200790
rect 311452 200086 311756 200114
rect 310888 197736 310940 197742
rect 310888 197678 310940 197684
rect 311728 5030 311756 200086
rect 311820 198558 311848 200790
rect 311808 198552 311860 198558
rect 311808 198494 311860 198500
rect 311992 198076 312044 198082
rect 311992 198018 312044 198024
rect 311808 197736 311860 197742
rect 311808 197678 311860 197684
rect 311820 5166 311848 197678
rect 312004 16574 312032 198018
rect 312372 197606 312400 200790
rect 312924 198694 312952 200790
rect 312912 198688 312964 198694
rect 312912 198630 312964 198636
rect 312544 198212 312596 198218
rect 312544 198154 312596 198160
rect 312360 197600 312412 197606
rect 312360 197542 312412 197548
rect 312004 16546 312216 16574
rect 311808 5160 311860 5166
rect 311808 5102 311860 5108
rect 311716 5024 311768 5030
rect 311716 4966 311768 4972
rect 311440 3392 311492 3398
rect 311440 3334 311492 3340
rect 310428 3324 310480 3330
rect 310428 3266 310480 3272
rect 310244 3188 310296 3194
rect 310244 3130 310296 3136
rect 310256 480 310284 3130
rect 311452 480 311480 3334
rect 312188 490 312216 16546
rect 312556 4146 312584 198154
rect 312544 4140 312596 4146
rect 312544 4082 312596 4088
rect 313200 3738 313228 200790
rect 314028 198014 314056 200790
rect 314016 198008 314068 198014
rect 314016 197950 314068 197956
rect 313924 197600 313976 197606
rect 313924 197542 313976 197548
rect 313936 5098 313964 197542
rect 313924 5092 313976 5098
rect 313924 5034 313976 5040
rect 314488 4894 314516 200790
rect 314568 198008 314620 198014
rect 314568 197950 314620 197956
rect 314580 4962 314608 197950
rect 314948 197470 314976 200790
rect 315500 197538 315528 200790
rect 315960 198286 315988 200790
rect 315948 198280 316000 198286
rect 315948 198222 316000 198228
rect 315488 197532 315540 197538
rect 315488 197474 315540 197480
rect 314936 197464 314988 197470
rect 314936 197406 314988 197412
rect 316604 197402 316632 200790
rect 317156 200114 317184 200790
rect 317156 200086 317276 200114
rect 316684 197464 316736 197470
rect 316684 197406 316736 197412
rect 316592 197396 316644 197402
rect 316592 197338 316644 197344
rect 314568 4956 314620 4962
rect 314568 4898 314620 4904
rect 314476 4888 314528 4894
rect 314476 4830 314528 4836
rect 316224 4140 316276 4146
rect 316224 4082 316276 4088
rect 313832 3936 313884 3942
rect 313832 3878 313884 3884
rect 313188 3732 313240 3738
rect 313188 3674 313240 3680
rect 312464 598 312676 626
rect 312464 490 312492 598
rect 298438 -960 298550 480
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301934 -960 302046 480
rect 303130 -960 303242 480
rect 304326 -960 304438 480
rect 305522 -960 305634 480
rect 306718 -960 306830 480
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 310214 -960 310326 480
rect 311410 -960 311522 480
rect 312188 462 312492 490
rect 312648 480 312676 598
rect 313844 480 313872 3878
rect 315028 3528 315080 3534
rect 315028 3470 315080 3476
rect 315040 480 315068 3470
rect 316236 480 316264 4082
rect 316696 3738 316724 197406
rect 317248 6186 317276 200086
rect 317340 198082 317368 200790
rect 317328 198076 317380 198082
rect 317328 198018 317380 198024
rect 317984 197402 318012 200790
rect 318536 198218 318564 200790
rect 319180 198626 319208 200790
rect 319168 198620 319220 198626
rect 319168 198562 319220 198568
rect 318524 198212 318576 198218
rect 318524 198154 318576 198160
rect 318064 198076 318116 198082
rect 318064 198018 318116 198024
rect 317328 197396 317380 197402
rect 317328 197338 317380 197344
rect 317972 197396 318024 197402
rect 317972 197338 318024 197344
rect 317236 6180 317288 6186
rect 317236 6122 317288 6128
rect 317340 5114 317368 197338
rect 317248 5086 317368 5114
rect 316684 3732 316736 3738
rect 316684 3674 316736 3680
rect 317248 3534 317276 5086
rect 318076 4826 318104 198018
rect 318156 197532 318208 197538
rect 318156 197474 318208 197480
rect 318168 14686 318196 197474
rect 319548 197402 319576 200790
rect 320100 198490 320128 200790
rect 320088 198484 320140 198490
rect 320088 198426 320140 198432
rect 320652 197742 320680 200790
rect 320640 197736 320692 197742
rect 320640 197678 320692 197684
rect 321112 197606 321140 200790
rect 321100 197600 321152 197606
rect 321100 197542 321152 197548
rect 318708 197396 318760 197402
rect 318708 197338 318760 197344
rect 319536 197396 319588 197402
rect 319536 197338 319588 197344
rect 318156 14680 318208 14686
rect 318156 14622 318208 14628
rect 318064 4820 318116 4826
rect 318064 4762 318116 4768
rect 318720 3806 318748 197338
rect 321296 14550 321324 200926
rect 321862 200790 322152 200818
rect 322414 200790 322796 200818
rect 322966 200790 323256 200818
rect 323426 200790 323808 200818
rect 323978 200790 324268 200818
rect 324530 200790 324912 200818
rect 324990 200790 325464 200818
rect 325542 200790 325648 200818
rect 326002 200790 326384 200818
rect 326554 200790 326936 200818
rect 327106 200790 327488 200818
rect 327566 200790 327856 200818
rect 328118 200790 328316 200818
rect 328578 200790 328960 200818
rect 329130 200790 329604 200818
rect 329682 200790 329788 200818
rect 330142 200790 330432 200818
rect 330694 200790 330984 200818
rect 331246 200790 331536 200818
rect 331706 200790 332088 200818
rect 332258 200790 332456 200818
rect 332718 200790 333008 200818
rect 333270 200790 333560 200818
rect 333822 200790 333928 200818
rect 334282 200790 334664 200818
rect 334834 200790 335032 200818
rect 322124 197878 322152 200790
rect 322112 197872 322164 197878
rect 322112 197814 322164 197820
rect 321468 197736 321520 197742
rect 321468 197678 321520 197684
rect 321376 197600 321428 197606
rect 321376 197542 321428 197548
rect 321284 14544 321336 14550
rect 321284 14486 321336 14492
rect 319720 4072 319772 4078
rect 319720 4014 319772 4020
rect 318524 3800 318576 3806
rect 318524 3742 318576 3748
rect 318708 3800 318760 3806
rect 318708 3742 318760 3748
rect 317236 3528 317288 3534
rect 317236 3470 317288 3476
rect 317328 3460 317380 3466
rect 317328 3402 317380 3408
rect 317340 480 317368 3402
rect 318536 480 318564 3742
rect 319732 480 319760 4014
rect 320916 4004 320968 4010
rect 320916 3946 320968 3952
rect 320928 480 320956 3946
rect 321388 3126 321416 197542
rect 321376 3120 321428 3126
rect 321376 3062 321428 3068
rect 321480 3058 321508 197678
rect 322204 197396 322256 197402
rect 322204 197338 322256 197344
rect 322112 3596 322164 3602
rect 322112 3538 322164 3544
rect 321468 3052 321520 3058
rect 321468 2994 321520 3000
rect 322124 480 322152 3538
rect 322216 2990 322244 197338
rect 322768 3602 322796 200790
rect 323124 198144 323176 198150
rect 323124 198086 323176 198092
rect 322848 197872 322900 197878
rect 322848 197814 322900 197820
rect 322756 3596 322808 3602
rect 322756 3538 322808 3544
rect 322860 3194 322888 197814
rect 323136 190454 323164 198086
rect 323228 197470 323256 200790
rect 323216 197464 323268 197470
rect 323216 197406 323268 197412
rect 323780 197402 323808 200790
rect 324240 197538 324268 200790
rect 324228 197532 324280 197538
rect 324228 197474 324280 197480
rect 324136 197464 324188 197470
rect 324136 197406 324188 197412
rect 323768 197396 323820 197402
rect 323768 197338 323820 197344
rect 323136 190426 323256 190454
rect 323228 16574 323256 190426
rect 323228 16546 323348 16574
rect 322848 3188 322900 3194
rect 322848 3130 322900 3136
rect 322204 2984 322256 2990
rect 322204 2926 322256 2932
rect 323320 480 323348 16546
rect 324148 14618 324176 197406
rect 324884 197402 324912 200790
rect 325436 197606 325464 200790
rect 325620 200114 325648 200790
rect 325528 200086 325648 200114
rect 325424 197600 325476 197606
rect 325424 197542 325476 197548
rect 324228 197396 324280 197402
rect 324228 197338 324280 197344
rect 324872 197396 324924 197402
rect 324872 197338 324924 197344
rect 325424 197396 325476 197402
rect 325424 197338 325476 197344
rect 324136 14612 324188 14618
rect 324136 14554 324188 14560
rect 324240 3398 324268 197338
rect 325436 11898 325464 197338
rect 325424 11892 325476 11898
rect 325424 11834 325476 11840
rect 325528 11778 325556 200086
rect 326356 197810 326384 200790
rect 326908 198354 326936 200790
rect 326896 198348 326948 198354
rect 326896 198290 326948 198296
rect 327460 198150 327488 200790
rect 327448 198144 327500 198150
rect 327448 198086 327500 198092
rect 327724 198008 327776 198014
rect 327724 197950 327776 197956
rect 326344 197804 326396 197810
rect 326344 197746 326396 197752
rect 325608 197600 325660 197606
rect 325608 197542 325660 197548
rect 325436 11750 325556 11778
rect 324412 5296 324464 5302
rect 324412 5238 324464 5244
rect 324228 3392 324280 3398
rect 324228 3334 324280 3340
rect 324424 480 324452 5238
rect 325436 3330 325464 11750
rect 325620 6914 325648 197542
rect 325528 6886 325648 6914
rect 325424 3324 325476 3330
rect 325424 3266 325476 3272
rect 325528 3262 325556 6886
rect 325608 3936 325660 3942
rect 325608 3878 325660 3884
rect 325516 3256 325568 3262
rect 325516 3198 325568 3204
rect 325620 480 325648 3878
rect 326804 3868 326856 3874
rect 326804 3810 326856 3816
rect 326816 480 326844 3810
rect 327736 3738 327764 197950
rect 327828 197402 327856 200790
rect 327908 198280 327960 198286
rect 327908 198222 327960 198228
rect 327816 197396 327868 197402
rect 327816 197338 327868 197344
rect 327920 180794 327948 198222
rect 328288 197742 328316 200790
rect 328932 197878 328960 200790
rect 329576 200114 329604 200790
rect 329576 200086 329696 200114
rect 328920 197872 328972 197878
rect 328920 197814 328972 197820
rect 328276 197736 328328 197742
rect 328276 197678 328328 197684
rect 328368 197396 328420 197402
rect 328368 197338 328420 197344
rect 327828 180766 327948 180794
rect 327828 5234 327856 180766
rect 328380 11762 328408 197338
rect 329668 14482 329696 200086
rect 329760 198014 329788 200790
rect 329748 198008 329800 198014
rect 329748 197950 329800 197956
rect 329748 197872 329800 197878
rect 329748 197814 329800 197820
rect 329656 14476 329708 14482
rect 329656 14418 329708 14424
rect 328368 11756 328420 11762
rect 328368 11698 328420 11704
rect 327816 5228 327868 5234
rect 327816 5170 327868 5176
rect 328000 5160 328052 5166
rect 328000 5102 328052 5108
rect 327724 3732 327776 3738
rect 327724 3674 327776 3680
rect 328012 480 328040 5102
rect 329760 4078 329788 197814
rect 330404 197402 330432 200790
rect 330484 198552 330536 198558
rect 330484 198494 330536 198500
rect 330392 197396 330444 197402
rect 330392 197338 330444 197344
rect 329748 4072 329800 4078
rect 329748 4014 329800 4020
rect 329196 3868 329248 3874
rect 329196 3810 329248 3816
rect 329208 480 329236 3810
rect 330496 3738 330524 198494
rect 330956 198286 330984 200790
rect 330944 198280 330996 198286
rect 330944 198222 330996 198228
rect 331508 197402 331536 200790
rect 332060 197470 332088 200790
rect 332048 197464 332100 197470
rect 332048 197406 332100 197412
rect 331128 197396 331180 197402
rect 331128 197338 331180 197344
rect 331496 197396 331548 197402
rect 331496 197338 331548 197344
rect 332324 197396 332376 197402
rect 332324 197338 332376 197344
rect 331140 4146 331168 197338
rect 331588 5092 331640 5098
rect 331588 5034 331640 5040
rect 331128 4140 331180 4146
rect 331128 4082 331180 4088
rect 330392 3732 330444 3738
rect 330392 3674 330444 3680
rect 330484 3732 330536 3738
rect 330484 3674 330536 3680
rect 330404 480 330432 3674
rect 331600 480 331628 5034
rect 332336 4350 332364 197338
rect 332428 4418 332456 200790
rect 332980 198558 333008 200790
rect 332968 198552 333020 198558
rect 332968 198494 333020 198500
rect 333532 197878 333560 200790
rect 333520 197872 333572 197878
rect 333520 197814 333572 197820
rect 332508 197464 332560 197470
rect 332508 197406 332560 197412
rect 332416 4412 332468 4418
rect 332416 4354 332468 4360
rect 332324 4344 332376 4350
rect 332324 4286 332376 4292
rect 332520 4010 332548 197406
rect 332692 5024 332744 5030
rect 332692 4966 332744 4972
rect 332508 4004 332560 4010
rect 332508 3946 332560 3952
rect 332704 480 332732 4966
rect 333900 4486 333928 200790
rect 334636 197470 334664 200790
rect 334624 197464 334676 197470
rect 334624 197406 334676 197412
rect 335004 197402 335032 200790
rect 334992 197396 335044 197402
rect 334992 197338 335044 197344
rect 334992 4752 335044 4758
rect 334992 4694 335044 4700
rect 333888 4480 333940 4486
rect 333888 4422 333940 4428
rect 333888 3732 333940 3738
rect 333888 3674 333940 3680
rect 333900 480 333928 3674
rect 335004 2530 335032 4694
rect 335096 4690 335124 200926
rect 335846 200790 336136 200818
rect 336398 200790 336688 200818
rect 336858 200790 337240 200818
rect 337410 200790 337792 200818
rect 337870 200790 337976 200818
rect 338422 200790 338712 200818
rect 338974 200790 339264 200818
rect 335544 198688 335596 198694
rect 335544 198630 335596 198636
rect 335176 197464 335228 197470
rect 335176 197406 335228 197412
rect 335084 4684 335136 4690
rect 335084 4626 335136 4632
rect 335188 4554 335216 197406
rect 335268 197396 335320 197402
rect 335268 197338 335320 197344
rect 335176 4548 335228 4554
rect 335176 4490 335228 4496
rect 335280 3942 335308 197338
rect 335556 16574 335584 198630
rect 336004 198620 336056 198626
rect 336004 198562 336056 198568
rect 335556 16546 335952 16574
rect 335268 3936 335320 3942
rect 335268 3878 335320 3884
rect 335924 2802 335952 16546
rect 336016 2922 336044 198562
rect 336108 197470 336136 200790
rect 336096 197464 336148 197470
rect 336096 197406 336148 197412
rect 336660 3874 336688 200790
rect 337212 197402 337240 200790
rect 337200 197396 337252 197402
rect 337200 197338 337252 197344
rect 337764 190454 337792 200790
rect 337948 198694 337976 200790
rect 337936 198688 337988 198694
rect 337936 198630 337988 198636
rect 338684 197402 338712 200790
rect 338764 198484 338816 198490
rect 338764 198426 338816 198432
rect 338028 197396 338080 197402
rect 338028 197338 338080 197344
rect 338672 197396 338724 197402
rect 338672 197338 338724 197344
rect 337764 190426 337976 190454
rect 337948 4758 337976 190426
rect 337936 4752 337988 4758
rect 337936 4694 337988 4700
rect 338040 4622 338068 197338
rect 338776 6322 338804 198426
rect 339236 197946 339264 200790
rect 339328 200114 339356 200926
rect 339986 200790 340460 200818
rect 340538 200790 340828 200818
rect 340998 200790 341288 200818
rect 341550 200790 341932 200818
rect 342010 200790 342208 200818
rect 342562 200790 342944 200818
rect 343114 200790 343312 200818
rect 340432 200114 340460 200790
rect 339328 200086 339448 200114
rect 340432 200086 340736 200114
rect 339224 197940 339276 197946
rect 339224 197882 339276 197888
rect 339316 197396 339368 197402
rect 339316 197338 339368 197344
rect 338764 6316 338816 6322
rect 338764 6258 338816 6264
rect 339328 5506 339356 197338
rect 339316 5500 339368 5506
rect 339316 5442 339368 5448
rect 338672 4956 338724 4962
rect 338672 4898 338724 4904
rect 338028 4616 338080 4622
rect 338028 4558 338080 4564
rect 336648 3868 336700 3874
rect 336648 3810 336700 3816
rect 337476 3664 337528 3670
rect 337476 3606 337528 3612
rect 336004 2916 336056 2922
rect 336004 2858 336056 2864
rect 335924 2774 336320 2802
rect 335004 2502 335124 2530
rect 335096 480 335124 2502
rect 336292 480 336320 2774
rect 337488 480 337516 3606
rect 338684 480 338712 4898
rect 339420 3670 339448 200086
rect 340236 198552 340288 198558
rect 340236 198494 340288 198500
rect 340144 197804 340196 197810
rect 340144 197746 340196 197752
rect 340156 6254 340184 197746
rect 340248 86290 340276 198494
rect 340236 86284 340288 86290
rect 340236 86226 340288 86232
rect 340144 6248 340196 6254
rect 340144 6190 340196 6196
rect 340708 5438 340736 200086
rect 340696 5432 340748 5438
rect 340696 5374 340748 5380
rect 340800 5370 340828 200790
rect 341260 197402 341288 200790
rect 341904 200114 341932 200790
rect 341904 200086 342116 200114
rect 341524 197736 341576 197742
rect 341524 197678 341576 197684
rect 341248 197396 341300 197402
rect 341248 197338 341300 197344
rect 341536 17270 341564 197678
rect 341616 197464 341668 197470
rect 341616 197406 341668 197412
rect 341628 86562 341656 197406
rect 341616 86556 341668 86562
rect 341616 86498 341668 86504
rect 341524 17264 341576 17270
rect 341524 17206 341576 17212
rect 341984 14680 342036 14686
rect 341984 14622 342036 14628
rect 340788 5364 340840 5370
rect 340788 5306 340840 5312
rect 339868 4888 339920 4894
rect 339868 4830 339920 4836
rect 339408 3664 339460 3670
rect 339408 3606 339460 3612
rect 339880 480 339908 4830
rect 340972 3528 341024 3534
rect 340972 3470 341024 3476
rect 341996 3482 342024 14622
rect 342088 5302 342116 200086
rect 342180 197810 342208 200790
rect 342168 197804 342220 197810
rect 342168 197746 342220 197752
rect 342916 197402 342944 200790
rect 343284 197742 343312 200790
rect 343272 197736 343324 197742
rect 343272 197678 343324 197684
rect 342168 197396 342220 197402
rect 342168 197338 342220 197344
rect 342904 197396 342956 197402
rect 342904 197338 342956 197344
rect 342076 5296 342128 5302
rect 342076 5238 342128 5244
rect 342180 3738 342208 197338
rect 343272 5228 343324 5234
rect 343272 5170 343324 5176
rect 342168 3732 342220 3738
rect 342168 3674 342220 3680
rect 340984 480 341012 3470
rect 341996 3454 342208 3482
rect 342180 480 342208 3454
rect 343284 2666 343312 5170
rect 343376 5030 343404 200926
rect 344126 200790 344416 200818
rect 344586 200790 344968 200818
rect 345138 200790 345520 200818
rect 345690 200790 346072 200818
rect 346150 200790 346256 200818
rect 346702 200790 346992 200818
rect 347254 200790 347544 200818
rect 344388 198422 344416 200790
rect 344376 198416 344428 198422
rect 344376 198358 344428 198364
rect 343456 197736 343508 197742
rect 343456 197678 343508 197684
rect 343468 5234 343496 197678
rect 343548 197396 343600 197402
rect 343548 197338 343600 197344
rect 343456 5228 343508 5234
rect 343456 5170 343508 5176
rect 343364 5024 343416 5030
rect 343364 4966 343416 4972
rect 343560 3534 343588 197338
rect 344940 5166 344968 200790
rect 345492 197470 345520 200790
rect 345480 197464 345532 197470
rect 345480 197406 345532 197412
rect 346044 197402 346072 200790
rect 346228 200114 346256 200790
rect 346136 200086 346256 200114
rect 346032 197396 346084 197402
rect 346032 197338 346084 197344
rect 345756 6180 345808 6186
rect 345756 6122 345808 6128
rect 344928 5160 344980 5166
rect 344928 5102 344980 5108
rect 343548 3528 343600 3534
rect 343548 3470 343600 3476
rect 344560 3460 344612 3466
rect 344560 3402 344612 3408
rect 343284 2638 343404 2666
rect 343376 480 343404 2638
rect 344572 480 344600 3402
rect 345768 480 345796 6122
rect 346136 4962 346164 200086
rect 346216 197464 346268 197470
rect 346216 197406 346268 197412
rect 346228 5098 346256 197406
rect 346964 197402 346992 200790
rect 347516 198626 347544 200790
rect 347608 200114 347636 200926
rect 348266 200790 348648 200818
rect 348726 200790 349016 200818
rect 349278 200790 349568 200818
rect 349830 200790 350212 200818
rect 350290 200790 350488 200818
rect 350842 200790 351224 200818
rect 351302 200790 351592 200818
rect 347608 200086 347728 200114
rect 347504 198620 347556 198626
rect 347504 198562 347556 198568
rect 346308 197396 346360 197402
rect 346308 197338 346360 197344
rect 346952 197396 347004 197402
rect 346952 197338 347004 197344
rect 347596 197396 347648 197402
rect 347596 197338 347648 197344
rect 346216 5092 346268 5098
rect 346216 5034 346268 5040
rect 346124 4956 346176 4962
rect 346124 4898 346176 4904
rect 346320 3466 346348 197338
rect 346952 4820 347004 4826
rect 346952 4762 347004 4768
rect 346308 3460 346360 3466
rect 346308 3402 346360 3408
rect 346964 480 346992 4762
rect 347608 4214 347636 197338
rect 347700 4894 347728 200086
rect 348620 197402 348648 200790
rect 348988 197742 349016 200790
rect 349344 198212 349396 198218
rect 349344 198154 349396 198160
rect 348976 197736 349028 197742
rect 348976 197678 349028 197684
rect 348608 197396 348660 197402
rect 348608 197338 348660 197344
rect 349068 197396 349120 197402
rect 349068 197338 349120 197344
rect 347688 4888 347740 4894
rect 347688 4830 347740 4836
rect 349080 4826 349108 197338
rect 349356 6914 349384 198154
rect 349540 197402 349568 200790
rect 350184 197554 350212 200790
rect 350460 198558 350488 200790
rect 350448 198552 350500 198558
rect 350448 198494 350500 198500
rect 350184 197526 350488 197554
rect 349528 197396 349580 197402
rect 349528 197338 349580 197344
rect 350356 197396 350408 197402
rect 350356 197338 350408 197344
rect 350368 9382 350396 197338
rect 350356 9376 350408 9382
rect 350356 9318 350408 9324
rect 350460 7070 350488 197526
rect 351196 197470 351224 200790
rect 351564 200114 351592 200790
rect 351748 200410 351776 200926
rect 352406 200790 352696 200818
rect 352866 200790 353248 200818
rect 353418 200790 353800 200818
rect 353878 200790 354352 200818
rect 354430 200790 354628 200818
rect 354982 200790 355272 200818
rect 355442 200790 355824 200818
rect 351748 200382 351868 200410
rect 351564 200086 351776 200114
rect 351184 197464 351236 197470
rect 351184 197406 351236 197412
rect 351748 190454 351776 200086
rect 351840 198218 351868 200382
rect 352564 198416 352616 198422
rect 352564 198358 352616 198364
rect 351828 198212 351880 198218
rect 351828 198154 351880 198160
rect 351748 190426 351868 190454
rect 351840 7138 351868 190426
rect 351828 7132 351880 7138
rect 351828 7074 351880 7080
rect 350448 7064 350500 7070
rect 350448 7006 350500 7012
rect 349264 6886 349384 6914
rect 349068 4820 349120 4826
rect 349068 4762 349120 4768
rect 347596 4208 347648 4214
rect 347596 4150 347648 4156
rect 348056 3800 348108 3806
rect 348056 3742 348108 3748
rect 348068 480 348096 3742
rect 349264 480 349292 6886
rect 352576 3806 352604 198358
rect 352668 197402 352696 200790
rect 352656 197396 352708 197402
rect 352656 197338 352708 197344
rect 353116 197396 353168 197402
rect 353116 197338 353168 197344
rect 353128 9314 353156 197338
rect 353116 9308 353168 9314
rect 353116 9250 353168 9256
rect 353220 7206 353248 200790
rect 353772 198490 353800 200790
rect 354324 200114 354352 200790
rect 354324 200086 354536 200114
rect 353760 198484 353812 198490
rect 353760 198426 353812 198432
rect 353944 198348 353996 198354
rect 353944 198290 353996 198296
rect 353208 7200 353260 7206
rect 353208 7142 353260 7148
rect 352840 6316 352892 6322
rect 352840 6258 352892 6264
rect 352564 3800 352616 3806
rect 352564 3742 352616 3748
rect 351644 2984 351696 2990
rect 351644 2926 351696 2932
rect 350448 2916 350500 2922
rect 350448 2858 350500 2864
rect 350460 480 350488 2858
rect 351656 480 351684 2926
rect 352852 480 352880 6258
rect 353956 2922 353984 198290
rect 354508 17338 354536 200086
rect 354496 17332 354548 17338
rect 354496 17274 354548 17280
rect 354600 7274 354628 200790
rect 355244 197402 355272 200790
rect 355796 198286 355824 200790
rect 355888 200114 355916 200926
rect 356546 200790 356928 200818
rect 357006 200790 357388 200818
rect 357558 200790 357848 200818
rect 358018 200790 358400 200818
rect 358570 200790 358768 200818
rect 359122 200790 359412 200818
rect 359582 200790 359872 200818
rect 355888 200086 356008 200114
rect 355784 198280 355836 198286
rect 355784 198222 355836 198228
rect 355232 197396 355284 197402
rect 355232 197338 355284 197344
rect 355980 7342 356008 200086
rect 356900 198422 356928 200790
rect 356888 198416 356940 198422
rect 356888 198358 356940 198364
rect 356704 197532 356756 197538
rect 356704 197474 356756 197480
rect 356336 14544 356388 14550
rect 356336 14486 356388 14492
rect 355968 7336 356020 7342
rect 355968 7278 356020 7284
rect 354588 7268 354640 7274
rect 354588 7210 354640 7216
rect 355232 3120 355284 3126
rect 355232 3062 355284 3068
rect 354036 3052 354088 3058
rect 354036 2994 354088 3000
rect 353944 2916 353996 2922
rect 353944 2858 353996 2864
rect 354048 480 354076 2994
rect 355244 480 355272 3062
rect 356348 480 356376 14486
rect 356716 3126 356744 197474
rect 356796 197464 356848 197470
rect 356796 197406 356848 197412
rect 356808 19990 356836 197406
rect 356796 19984 356848 19990
rect 356796 19926 356848 19932
rect 357360 14822 357388 200790
rect 357820 198082 357848 200790
rect 358176 198280 358228 198286
rect 358176 198222 358228 198228
rect 357808 198076 357860 198082
rect 357808 198018 357860 198024
rect 358084 197736 358136 197742
rect 358084 197678 358136 197684
rect 357348 14816 357400 14822
rect 357348 14758 357400 14764
rect 358096 6914 358124 197678
rect 358188 10470 358216 198222
rect 358372 197674 358400 200790
rect 358360 197668 358412 197674
rect 358360 197610 358412 197616
rect 358268 14612 358320 14618
rect 358268 14554 358320 14560
rect 358176 10464 358228 10470
rect 358176 10406 358228 10412
rect 358096 6886 358216 6914
rect 357716 3596 357768 3602
rect 357716 3538 357768 3544
rect 357532 3188 357584 3194
rect 357532 3130 357584 3136
rect 356704 3120 356756 3126
rect 356704 3062 356756 3068
rect 357544 480 357572 3130
rect 357728 2854 357756 3538
rect 358188 3194 358216 6886
rect 358280 3602 358308 14554
rect 358740 13122 358768 200790
rect 358820 198144 358872 198150
rect 358820 198086 358872 198092
rect 358832 197538 358860 198086
rect 359384 197742 359412 200790
rect 359844 198354 359872 200790
rect 360028 200114 360056 200926
rect 360594 200790 360976 200818
rect 361146 200790 361528 200818
rect 361698 200790 362080 200818
rect 362158 200790 362448 200818
rect 362710 200790 362908 200818
rect 363262 200790 363552 200818
rect 363722 200790 364104 200818
rect 360028 200086 360148 200114
rect 359832 198348 359884 198354
rect 359832 198290 359884 198296
rect 359464 198212 359516 198218
rect 359464 198154 359516 198160
rect 359372 197736 359424 197742
rect 359372 197678 359424 197684
rect 358820 197532 358872 197538
rect 358820 197474 358872 197480
rect 358728 13116 358780 13122
rect 358728 13058 358780 13064
rect 358268 3596 358320 3602
rect 358268 3538 358320 3544
rect 358176 3188 358228 3194
rect 358176 3130 358228 3136
rect 359476 2990 359504 198154
rect 359556 197532 359608 197538
rect 359556 197474 359608 197480
rect 359464 2984 359516 2990
rect 359464 2926 359516 2932
rect 359568 2854 359596 197474
rect 360120 9178 360148 200086
rect 360948 198014 360976 200790
rect 361028 198280 361080 198286
rect 361028 198222 361080 198228
rect 360936 198008 360988 198014
rect 360936 197950 360988 197956
rect 360936 197872 360988 197878
rect 360936 197814 360988 197820
rect 360844 197396 360896 197402
rect 360844 197338 360896 197344
rect 360108 9172 360160 9178
rect 360108 9114 360160 9120
rect 359924 3596 359976 3602
rect 359924 3538 359976 3544
rect 357716 2848 357768 2854
rect 357716 2790 357768 2796
rect 358728 2848 358780 2854
rect 358728 2790 358780 2796
rect 359556 2848 359608 2854
rect 359556 2790 359608 2796
rect 358740 480 358768 2790
rect 359936 480 359964 3538
rect 360856 3058 360884 197338
rect 360948 3194 360976 197814
rect 361040 14550 361068 198222
rect 361500 197470 361528 200790
rect 361488 197464 361540 197470
rect 361488 197406 361540 197412
rect 362052 197402 362080 200790
rect 362420 197538 362448 200790
rect 362880 198286 362908 200790
rect 362868 198280 362920 198286
rect 362868 198222 362920 198228
rect 362408 197532 362460 197538
rect 362408 197474 362460 197480
rect 363524 197402 363552 200790
rect 363696 198144 363748 198150
rect 363696 198086 363748 198092
rect 363604 197464 363656 197470
rect 363604 197406 363656 197412
rect 362040 197396 362092 197402
rect 362040 197338 362092 197344
rect 362868 197396 362920 197402
rect 362868 197338 362920 197344
rect 363512 197396 363564 197402
rect 363512 197338 363564 197344
rect 362880 86426 362908 197338
rect 362868 86420 362920 86426
rect 362868 86362 362920 86368
rect 361028 14544 361080 14550
rect 361028 14486 361080 14492
rect 363512 11824 363564 11830
rect 363512 11766 363564 11772
rect 361120 3392 361172 3398
rect 361120 3334 361172 3340
rect 360936 3188 360988 3194
rect 360936 3130 360988 3136
rect 360844 3052 360896 3058
rect 360844 2994 360896 3000
rect 361132 480 361160 3334
rect 362316 3120 362368 3126
rect 362316 3062 362368 3068
rect 362328 480 362356 3062
rect 363524 480 363552 11766
rect 363616 3398 363644 197406
rect 363708 10334 363736 198086
rect 364076 197470 364104 200790
rect 364168 197606 364196 200926
rect 364734 200790 365024 200818
rect 365286 200790 365576 200818
rect 365838 200790 366128 200818
rect 366298 200790 366772 200818
rect 366850 200790 366956 200818
rect 367310 200790 367600 200818
rect 367862 200790 368152 200818
rect 364892 197668 364944 197674
rect 364892 197610 364944 197616
rect 364156 197600 364208 197606
rect 364156 197542 364208 197548
rect 364064 197464 364116 197470
rect 364064 197406 364116 197412
rect 364248 197396 364300 197402
rect 364248 197338 364300 197344
rect 363696 10328 363748 10334
rect 363696 10270 363748 10276
rect 364260 5642 364288 197338
rect 364904 190454 364932 197610
rect 364996 197402 365024 200790
rect 365548 197674 365576 200790
rect 366100 198082 366128 200790
rect 366088 198076 366140 198082
rect 366088 198018 366140 198024
rect 365536 197668 365588 197674
rect 365536 197610 365588 197616
rect 366364 197532 366416 197538
rect 366364 197474 366416 197480
rect 364984 197396 365036 197402
rect 364984 197338 365036 197344
rect 365628 197396 365680 197402
rect 365628 197338 365680 197344
rect 364904 190426 365024 190454
rect 364248 5636 364300 5642
rect 364248 5578 364300 5584
rect 363604 3392 363656 3398
rect 363604 3334 363656 3340
rect 364616 3256 364668 3262
rect 364616 3198 364668 3204
rect 364628 480 364656 3198
rect 364996 3194 365024 190426
rect 365640 5710 365668 197338
rect 366376 86494 366404 197474
rect 366744 190454 366772 200790
rect 366928 198218 366956 200790
rect 366916 198212 366968 198218
rect 366916 198154 366968 198160
rect 367572 197878 367600 200790
rect 368124 200114 368152 200790
rect 368308 200410 368336 200926
rect 368874 200790 369256 200818
rect 369426 200790 369808 200818
rect 369886 200790 370176 200818
rect 370438 200790 370912 200818
rect 370990 200790 371188 200818
rect 371450 200790 371832 200818
rect 372002 200790 372384 200818
rect 368308 200382 368428 200410
rect 368124 200086 368336 200114
rect 367744 197940 367796 197946
rect 367744 197882 367796 197888
rect 367560 197872 367612 197878
rect 367560 197814 367612 197820
rect 366744 190426 367048 190454
rect 366364 86488 366416 86494
rect 366364 86430 366416 86436
rect 366916 6248 366968 6254
rect 366916 6190 366968 6196
rect 365628 5704 365680 5710
rect 365628 5646 365680 5652
rect 365812 3324 365864 3330
rect 365812 3266 365864 3272
rect 364984 3188 365036 3194
rect 364984 3130 365036 3136
rect 365824 480 365852 3266
rect 366928 3210 366956 6190
rect 367020 5778 367048 190426
rect 367756 6186 367784 197882
rect 367836 197804 367888 197810
rect 367836 197746 367888 197752
rect 367848 10402 367876 197746
rect 368308 190454 368336 200086
rect 368400 197402 368428 200382
rect 369228 197946 369256 200790
rect 369216 197940 369268 197946
rect 369216 197882 369268 197888
rect 368388 197396 368440 197402
rect 368388 197338 368440 197344
rect 368308 190426 368428 190454
rect 367928 14476 367980 14482
rect 367928 14418 367980 14424
rect 367836 10396 367888 10402
rect 367836 10338 367888 10344
rect 367744 6180 367796 6186
rect 367744 6122 367796 6128
rect 367008 5772 367060 5778
rect 367008 5714 367060 5720
rect 367940 4282 367968 14418
rect 368400 5846 368428 190426
rect 369780 5914 369808 200790
rect 370148 197878 370176 200790
rect 370596 198144 370648 198150
rect 370596 198086 370648 198092
rect 370136 197872 370188 197878
rect 370136 197814 370188 197820
rect 370504 197396 370556 197402
rect 370504 197338 370556 197344
rect 370516 25566 370544 197338
rect 370608 35222 370636 198086
rect 370884 198082 370912 200790
rect 370872 198076 370924 198082
rect 370872 198018 370924 198024
rect 370688 197464 370740 197470
rect 370688 197406 370740 197412
rect 370700 84930 370728 197406
rect 370688 84924 370740 84930
rect 370688 84866 370740 84872
rect 370596 35216 370648 35222
rect 370596 35158 370648 35164
rect 370504 25560 370556 25566
rect 370504 25502 370556 25508
rect 370136 11756 370188 11762
rect 370136 11698 370188 11704
rect 369768 5908 369820 5914
rect 369768 5850 369820 5856
rect 368388 5840 368440 5846
rect 368388 5782 368440 5788
rect 367928 4276 367980 4282
rect 367928 4218 367980 4224
rect 366928 3182 367048 3210
rect 367020 480 367048 3182
rect 368204 2916 368256 2922
rect 368204 2858 368256 2864
rect 368216 480 368244 2858
rect 369400 2848 369452 2854
rect 369400 2790 369452 2796
rect 369412 480 369440 2790
rect 370148 490 370176 11698
rect 371160 5982 371188 200790
rect 371804 197538 371832 200790
rect 371976 198008 372028 198014
rect 371976 197950 372028 197956
rect 371884 197736 371936 197742
rect 371884 197678 371936 197684
rect 371792 197532 371844 197538
rect 371792 197474 371844 197480
rect 371240 17264 371292 17270
rect 371240 17206 371292 17212
rect 371148 5976 371200 5982
rect 371148 5918 371200 5924
rect 370424 598 370636 626
rect 370424 490 370452 598
rect 312606 -960 312718 480
rect 313802 -960 313914 480
rect 314998 -960 315110 480
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318494 -960 318606 480
rect 319690 -960 319802 480
rect 320886 -960 320998 480
rect 322082 -960 322194 480
rect 323278 -960 323390 480
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326774 -960 326886 480
rect 327970 -960 328082 480
rect 329166 -960 329278 480
rect 330362 -960 330474 480
rect 331558 -960 331670 480
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 335054 -960 335166 480
rect 336250 -960 336362 480
rect 337446 -960 337558 480
rect 338642 -960 338754 480
rect 339838 -960 339950 480
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 343334 -960 343446 480
rect 344530 -960 344642 480
rect 345726 -960 345838 480
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351614 -960 351726 480
rect 352810 -960 352922 480
rect 354006 -960 354118 480
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359894 -960 360006 480
rect 361090 -960 361202 480
rect 362286 -960 362398 480
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 368174 -960 368286 480
rect 369370 -960 369482 480
rect 370148 462 370452 490
rect 370608 480 370636 598
rect 371252 490 371280 17206
rect 371896 16182 371924 197678
rect 371884 16176 371936 16182
rect 371884 16118 371936 16124
rect 371988 16114 372016 197950
rect 372356 197674 372384 200790
rect 372448 200114 372476 200926
rect 373014 200790 373304 200818
rect 373566 200790 373856 200818
rect 374026 200790 374408 200818
rect 374578 200790 374960 200818
rect 375130 200790 375328 200818
rect 375590 200790 375880 200818
rect 376142 200790 376524 200818
rect 376602 200790 376708 200818
rect 377154 200790 377536 200818
rect 377706 200790 378088 200818
rect 378166 200790 378456 200818
rect 378718 200790 379100 200818
rect 379178 200790 379468 200818
rect 379730 200790 380112 200818
rect 380282 200790 380664 200818
rect 380742 200790 380848 200818
rect 381294 200790 381584 200818
rect 381846 200790 382228 200818
rect 382306 200790 382688 200818
rect 382858 200790 383240 200818
rect 383318 200790 383516 200818
rect 383870 200790 384160 200818
rect 384422 200790 384712 200818
rect 384882 200790 384988 200818
rect 385434 200790 385816 200818
rect 385894 200790 386184 200818
rect 386446 200790 386736 200818
rect 386998 200790 387380 200818
rect 387458 200790 387748 200818
rect 388010 200790 388392 200818
rect 388562 200790 388944 200818
rect 389022 200790 389128 200818
rect 389574 200790 389864 200818
rect 390034 200790 390416 200818
rect 390586 200790 390968 200818
rect 391138 200790 391520 200818
rect 391598 200790 391888 200818
rect 392150 200790 392440 200818
rect 392610 200790 393084 200818
rect 393162 200790 393268 200818
rect 393714 200790 394096 200818
rect 394174 200790 394648 200818
rect 394726 200790 395016 200818
rect 395186 200790 395568 200818
rect 395738 200790 396028 200818
rect 396290 200790 396672 200818
rect 396750 200790 397040 200818
rect 397302 200790 397408 200818
rect 397854 200790 398144 200818
rect 398314 200790 398696 200818
rect 398866 200790 399248 200818
rect 399326 200790 399616 200818
rect 399878 200790 400168 200818
rect 400430 200790 400720 200818
rect 400890 200790 401364 200818
rect 401442 200790 401548 200818
rect 401902 200790 402192 200818
rect 402454 200790 402836 200818
rect 403006 200790 403296 200818
rect 403466 200790 403848 200818
rect 404018 200790 404216 200818
rect 404570 200790 404952 200818
rect 405030 200790 405504 200818
rect 405582 200790 405688 200818
rect 406042 200790 406516 200818
rect 406594 200790 407068 200818
rect 407146 200790 407528 200818
rect 407606 200790 407896 200818
rect 408158 200790 408448 200818
rect 408618 200790 409000 200818
rect 409170 200790 409552 200818
rect 409722 200790 409828 200818
rect 410182 200790 410472 200818
rect 410734 200790 410932 200818
rect 372448 200086 372568 200114
rect 372068 197668 372120 197674
rect 372068 197610 372120 197616
rect 372344 197668 372396 197674
rect 372344 197610 372396 197616
rect 372080 87650 372108 197610
rect 372068 87644 372120 87650
rect 372068 87586 372120 87592
rect 371976 16108 372028 16114
rect 371976 16050 372028 16056
rect 372540 6118 372568 200086
rect 373276 197470 373304 200790
rect 373828 198014 373856 200790
rect 373816 198008 373868 198014
rect 373816 197950 373868 197956
rect 373264 197464 373316 197470
rect 373264 197406 373316 197412
rect 374380 197402 374408 200790
rect 374932 197470 374960 200790
rect 374644 197464 374696 197470
rect 374644 197406 374696 197412
rect 374920 197464 374972 197470
rect 374920 197406 374972 197412
rect 374368 197396 374420 197402
rect 374368 197338 374420 197344
rect 374656 10266 374684 197406
rect 375196 197396 375248 197402
rect 375196 197338 375248 197344
rect 375104 10328 375156 10334
rect 375104 10270 375156 10276
rect 374644 10260 374696 10266
rect 374644 10202 374696 10208
rect 372528 6112 372580 6118
rect 372528 6054 372580 6060
rect 374092 4140 374144 4146
rect 374092 4082 374144 4088
rect 372896 4072 372948 4078
rect 372896 4014 372948 4020
rect 371528 598 371740 626
rect 371528 490 371556 598
rect 370566 -960 370678 480
rect 371252 462 371556 490
rect 371712 480 371740 598
rect 372908 480 372936 4014
rect 374104 480 374132 4082
rect 375116 3482 375144 10270
rect 375208 6050 375236 197338
rect 375196 6044 375248 6050
rect 375196 5986 375248 5992
rect 375300 4078 375328 200790
rect 375852 197402 375880 200790
rect 376024 197600 376076 197606
rect 376024 197542 376076 197548
rect 375840 197396 375892 197402
rect 375840 197338 375892 197344
rect 375288 4072 375340 4078
rect 375288 4014 375340 4020
rect 375116 3454 375328 3482
rect 375300 480 375328 3454
rect 376036 3262 376064 197542
rect 376392 197396 376444 197402
rect 376392 197338 376444 197344
rect 376404 190454 376432 197338
rect 376496 195242 376524 200790
rect 376680 197742 376708 200790
rect 376668 197736 376720 197742
rect 376668 197678 376720 197684
rect 377404 197464 377456 197470
rect 377404 197406 377456 197412
rect 376496 195214 376708 195242
rect 376404 190426 376616 190454
rect 376588 9042 376616 190426
rect 376576 9036 376628 9042
rect 376576 8978 376628 8984
rect 376680 6798 376708 195214
rect 377416 9110 377444 197406
rect 377508 197402 377536 200790
rect 377496 197396 377548 197402
rect 377496 197338 377548 197344
rect 377956 197396 378008 197402
rect 377956 197338 378008 197344
rect 377968 16046 377996 197338
rect 377956 16040 378008 16046
rect 377956 15982 378008 15988
rect 377680 14544 377732 14550
rect 377680 14486 377732 14492
rect 377404 9104 377456 9110
rect 377404 9046 377456 9052
rect 376668 6792 376720 6798
rect 376668 6734 376720 6740
rect 376484 3324 376536 3330
rect 376484 3266 376536 3272
rect 376024 3256 376076 3262
rect 376024 3198 376076 3204
rect 376496 480 376524 3266
rect 377692 480 377720 14486
rect 378060 6730 378088 200790
rect 378428 197402 378456 200790
rect 379072 200114 379100 200790
rect 379072 200086 379376 200114
rect 378784 197804 378836 197810
rect 378784 197746 378836 197752
rect 378416 197396 378468 197402
rect 378416 197338 378468 197344
rect 378048 6724 378100 6730
rect 378048 6666 378100 6672
rect 378796 3330 378824 197746
rect 379244 197396 379296 197402
rect 379244 197338 379296 197344
rect 379256 86358 379284 197338
rect 379244 86352 379296 86358
rect 379244 86294 379296 86300
rect 379348 11830 379376 200086
rect 379336 11824 379388 11830
rect 379336 11766 379388 11772
rect 379440 6662 379468 200790
rect 380084 197742 380112 200790
rect 380072 197736 380124 197742
rect 380072 197678 380124 197684
rect 380636 196790 380664 200790
rect 380624 196784 380676 196790
rect 380624 196726 380676 196732
rect 380820 180794 380848 200790
rect 381452 197668 381504 197674
rect 381452 197610 381504 197616
rect 381464 190454 381492 197610
rect 381556 197402 381584 200790
rect 381544 197396 381596 197402
rect 381544 197338 381596 197344
rect 382096 197396 382148 197402
rect 382096 197338 382148 197344
rect 381464 190426 381584 190454
rect 380728 180766 380848 180794
rect 379428 6656 379480 6662
rect 379428 6598 379480 6604
rect 380728 6594 380756 180766
rect 380716 6588 380768 6594
rect 380716 6530 380768 6536
rect 381176 4412 381228 4418
rect 381176 4354 381228 4360
rect 378876 4344 378928 4350
rect 378876 4286 378928 4292
rect 378784 3324 378836 3330
rect 378784 3266 378836 3272
rect 378888 480 378916 4286
rect 379980 4004 380032 4010
rect 379980 3946 380032 3952
rect 379992 480 380020 3946
rect 381188 480 381216 4354
rect 381556 4146 381584 190426
rect 382108 21418 382136 197338
rect 382096 21412 382148 21418
rect 382096 21354 382148 21360
rect 382200 11762 382228 200790
rect 382660 197402 382688 200790
rect 383212 197674 383240 200790
rect 383200 197668 383252 197674
rect 383200 197610 383252 197616
rect 382648 197396 382700 197402
rect 382648 197338 382700 197344
rect 382372 86284 382424 86290
rect 382372 86226 382424 86232
rect 382188 11756 382240 11762
rect 382188 11698 382240 11704
rect 381544 4140 381596 4146
rect 381544 4082 381596 4088
rect 382384 480 382412 86226
rect 383488 8974 383516 200790
rect 384132 197402 384160 200790
rect 384684 197606 384712 200790
rect 384960 200114 384988 200790
rect 384868 200086 384988 200114
rect 384672 197600 384724 197606
rect 384672 197542 384724 197548
rect 383568 197396 383620 197402
rect 383568 197338 383620 197344
rect 384120 197396 384172 197402
rect 384120 197338 384172 197344
rect 383476 8968 383528 8974
rect 383476 8910 383528 8916
rect 383580 6526 383608 197338
rect 384868 89010 384896 200086
rect 385592 198212 385644 198218
rect 385592 198154 385644 198160
rect 384948 197396 385000 197402
rect 384948 197338 385000 197344
rect 384856 89004 384908 89010
rect 384856 88946 384908 88952
rect 383568 6520 383620 6526
rect 383568 6462 383620 6468
rect 384960 6458 384988 197338
rect 385604 190454 385632 198154
rect 385684 197532 385736 197538
rect 385684 197474 385736 197480
rect 385696 197282 385724 197474
rect 385788 197402 385816 200790
rect 386156 197538 386184 200790
rect 386144 197532 386196 197538
rect 386144 197474 386196 197480
rect 385776 197396 385828 197402
rect 385776 197338 385828 197344
rect 386328 197396 386380 197402
rect 386328 197338 386380 197344
rect 385696 197254 385816 197282
rect 385604 190426 385724 190454
rect 385696 9246 385724 190426
rect 385788 44878 385816 197254
rect 385776 44872 385828 44878
rect 385776 44814 385828 44820
rect 385684 9240 385736 9246
rect 385684 9182 385736 9188
rect 384948 6452 385000 6458
rect 384948 6394 385000 6400
rect 386340 6390 386368 197338
rect 386708 196722 386736 200790
rect 387352 200114 387380 200790
rect 387352 200086 387656 200114
rect 386696 196716 386748 196722
rect 386696 196658 386748 196664
rect 386328 6384 386380 6390
rect 386328 6326 386380 6332
rect 387628 6322 387656 200086
rect 387720 197470 387748 200790
rect 387708 197464 387760 197470
rect 387708 197406 387760 197412
rect 388364 197402 388392 200790
rect 388444 197600 388496 197606
rect 388444 197542 388496 197548
rect 388352 197396 388404 197402
rect 388352 197338 388404 197344
rect 388456 26926 388484 197542
rect 388536 197464 388588 197470
rect 388536 197406 388588 197412
rect 388548 86290 388576 197406
rect 388812 197396 388864 197402
rect 388812 197338 388864 197344
rect 388824 190454 388852 197338
rect 388916 195242 388944 200790
rect 389100 197538 389128 200790
rect 389088 197532 389140 197538
rect 389088 197474 389140 197480
rect 389836 197470 389864 200790
rect 389824 197464 389876 197470
rect 389824 197406 389876 197412
rect 388916 195214 389128 195242
rect 388824 190426 389036 190454
rect 388536 86284 388588 86290
rect 388536 86226 388588 86232
rect 388444 26920 388496 26926
rect 388444 26862 388496 26868
rect 389008 15910 389036 190426
rect 388996 15904 389048 15910
rect 388996 15846 389048 15852
rect 387616 6316 387668 6322
rect 387616 6258 387668 6264
rect 389100 6254 389128 195214
rect 389180 86556 389232 86562
rect 389180 86498 389232 86504
rect 389192 16574 389220 86498
rect 389192 16546 389496 16574
rect 389088 6248 389140 6254
rect 389088 6190 389140 6196
rect 388260 4684 388312 4690
rect 388260 4626 388312 4632
rect 385960 4548 386012 4554
rect 385960 4490 386012 4496
rect 384764 4480 384816 4486
rect 384764 4422 384816 4428
rect 383568 3120 383620 3126
rect 383568 3062 383620 3068
rect 383580 480 383608 3062
rect 384776 480 384804 4422
rect 385972 480 386000 4490
rect 387156 3936 387208 3942
rect 387156 3878 387208 3884
rect 387168 480 387196 3878
rect 388272 480 388300 4626
rect 389468 480 389496 16546
rect 390388 14618 390416 200790
rect 390468 197464 390520 197470
rect 390468 197406 390520 197412
rect 390376 14612 390428 14618
rect 390376 14554 390428 14560
rect 390480 4282 390508 197406
rect 390940 197402 390968 200790
rect 391492 200114 391520 200790
rect 391492 200086 391796 200114
rect 390928 197396 390980 197402
rect 390928 197338 390980 197344
rect 391768 4350 391796 200086
rect 391860 196654 391888 200790
rect 392412 198218 392440 200790
rect 392400 198212 392452 198218
rect 392400 198154 392452 198160
rect 393056 197402 393084 200790
rect 393240 200114 393268 200790
rect 393148 200086 393268 200114
rect 392584 197396 392636 197402
rect 392584 197338 392636 197344
rect 393044 197396 393096 197402
rect 393044 197338 393096 197344
rect 391848 196648 391900 196654
rect 391848 196590 391900 196596
rect 392596 24138 392624 197338
rect 392584 24132 392636 24138
rect 392584 24074 392636 24080
rect 393148 14482 393176 200086
rect 393504 198688 393556 198694
rect 393504 198630 393556 198636
rect 393228 197396 393280 197402
rect 393228 197338 393280 197344
rect 393136 14476 393188 14482
rect 393136 14418 393188 14424
rect 393044 4752 393096 4758
rect 393044 4694 393096 4700
rect 391848 4616 391900 4622
rect 391848 4558 391900 4564
rect 391756 4344 391808 4350
rect 391756 4286 391808 4292
rect 390468 4276 390520 4282
rect 390468 4218 390520 4224
rect 390652 3868 390704 3874
rect 390652 3810 390704 3816
rect 390664 480 390692 3810
rect 391860 480 391888 4558
rect 393056 480 393084 4694
rect 393240 4418 393268 197338
rect 393516 16574 393544 198630
rect 393964 197940 394016 197946
rect 393964 197882 394016 197888
rect 393516 16546 393912 16574
rect 393228 4412 393280 4418
rect 393228 4354 393280 4360
rect 393884 2938 393912 16546
rect 393976 3126 394004 197882
rect 394068 197402 394096 200790
rect 394056 197396 394108 197402
rect 394056 197338 394108 197344
rect 394620 4486 394648 200790
rect 394988 197878 395016 200790
rect 395540 198694 395568 200790
rect 395528 198688 395580 198694
rect 395528 198630 395580 198636
rect 394976 197872 395028 197878
rect 394976 197814 395028 197820
rect 395896 197872 395948 197878
rect 395896 197814 395948 197820
rect 395344 197396 395396 197402
rect 395344 197338 395396 197344
rect 395356 22778 395384 197338
rect 395344 22772 395396 22778
rect 395344 22714 395396 22720
rect 395908 14550 395936 197814
rect 395896 14544 395948 14550
rect 395896 14486 395948 14492
rect 395344 5500 395396 5506
rect 395344 5442 395396 5448
rect 394608 4480 394660 4486
rect 394608 4422 394660 4428
rect 393964 3120 394016 3126
rect 393964 3062 394016 3068
rect 393884 2910 394280 2938
rect 394252 480 394280 2910
rect 395356 480 395384 5442
rect 396000 4554 396028 200790
rect 396644 197402 396672 200790
rect 397012 197878 397040 200790
rect 397000 197872 397052 197878
rect 397000 197814 397052 197820
rect 396724 197600 396776 197606
rect 396724 197542 396776 197548
rect 396632 197396 396684 197402
rect 396632 197338 396684 197344
rect 396736 16250 396764 197542
rect 397276 197396 397328 197402
rect 397276 197338 397328 197344
rect 396724 16244 396776 16250
rect 396724 16186 396776 16192
rect 397288 7410 397316 197338
rect 397276 7404 397328 7410
rect 397276 7346 397328 7352
rect 396540 6180 396592 6186
rect 396540 6122 396592 6128
rect 395988 4548 396040 4554
rect 395988 4490 396040 4496
rect 396552 480 396580 6122
rect 397380 4622 397408 200790
rect 398116 197402 398144 200790
rect 398668 197538 398696 200790
rect 399220 197606 399248 200790
rect 399208 197600 399260 197606
rect 399208 197542 399260 197548
rect 398656 197532 398708 197538
rect 398656 197474 398708 197480
rect 399484 197532 399536 197538
rect 399484 197474 399536 197480
rect 398104 197396 398156 197402
rect 398104 197338 398156 197344
rect 398748 197396 398800 197402
rect 398748 197338 398800 197344
rect 398760 7478 398788 197338
rect 398748 7472 398800 7478
rect 398748 7414 398800 7420
rect 398932 5432 398984 5438
rect 398932 5374 398984 5380
rect 397368 4616 397420 4622
rect 397368 4558 397420 4564
rect 397736 3664 397788 3670
rect 397736 3606 397788 3612
rect 397748 480 397776 3606
rect 398944 480 398972 5374
rect 399496 4010 399524 197474
rect 399588 197402 399616 200790
rect 400140 198694 400168 200790
rect 400128 198688 400180 198694
rect 400128 198630 400180 198636
rect 400128 197600 400180 197606
rect 400128 197542 400180 197548
rect 399576 197396 399628 197402
rect 399576 197338 399628 197344
rect 400036 197396 400088 197402
rect 400036 197338 400088 197344
rect 400048 7546 400076 197338
rect 400036 7540 400088 7546
rect 400036 7482 400088 7488
rect 400140 6914 400168 197542
rect 400692 197402 400720 200790
rect 400864 197804 400916 197810
rect 400864 197746 400916 197752
rect 400680 197396 400732 197402
rect 400680 197338 400732 197344
rect 400876 84862 400904 197746
rect 400864 84856 400916 84862
rect 400864 84798 400916 84804
rect 401336 8294 401364 200790
rect 401416 197396 401468 197402
rect 401416 197338 401468 197344
rect 401324 8288 401376 8294
rect 401324 8230 401376 8236
rect 400048 6886 400168 6914
rect 400048 4690 400076 6886
rect 400128 5364 400180 5370
rect 400128 5306 400180 5312
rect 400036 4684 400088 4690
rect 400036 4626 400088 4632
rect 399484 4004 399536 4010
rect 399484 3946 399536 3952
rect 400140 480 400168 5306
rect 401428 4758 401456 197338
rect 401416 4752 401468 4758
rect 401416 4694 401468 4700
rect 401520 3942 401548 200790
rect 402164 197538 402192 200790
rect 402152 197532 402204 197538
rect 402152 197474 402204 197480
rect 402808 8226 402836 200790
rect 403268 197878 403296 200790
rect 403624 197940 403676 197946
rect 403624 197882 403676 197888
rect 403256 197872 403308 197878
rect 403256 197814 403308 197820
rect 402888 197532 402940 197538
rect 402888 197474 402940 197480
rect 402796 8220 402848 8226
rect 402796 8162 402848 8168
rect 402900 5506 402928 197474
rect 403636 16574 403664 197882
rect 403820 197538 403848 200790
rect 403808 197532 403860 197538
rect 403808 197474 403860 197480
rect 403636 16546 403756 16574
rect 403728 10402 403756 16546
rect 403624 10396 403676 10402
rect 403624 10338 403676 10344
rect 403716 10396 403768 10402
rect 403716 10338 403768 10344
rect 402888 5500 402940 5506
rect 402888 5442 402940 5448
rect 402520 5296 402572 5302
rect 402520 5238 402572 5244
rect 401508 3936 401560 3942
rect 401508 3878 401560 3884
rect 401324 3732 401376 3738
rect 401324 3674 401376 3680
rect 401336 480 401364 3674
rect 402532 480 402560 5238
rect 403636 480 403664 10338
rect 404188 8158 404216 200790
rect 404924 197538 404952 200790
rect 405476 197742 405504 200790
rect 405660 200114 405688 200790
rect 405568 200086 405688 200114
rect 406488 200114 406516 200790
rect 406488 200086 406608 200114
rect 405464 197736 405516 197742
rect 405464 197678 405516 197684
rect 404268 197532 404320 197538
rect 404268 197474 404320 197480
rect 404912 197532 404964 197538
rect 404912 197474 404964 197480
rect 404176 8152 404228 8158
rect 404176 8094 404228 8100
rect 404280 5438 404308 197474
rect 405568 8090 405596 200086
rect 405648 197736 405700 197742
rect 405648 197678 405700 197684
rect 405556 8084 405608 8090
rect 405556 8026 405608 8032
rect 404268 5432 404320 5438
rect 404268 5374 404320 5380
rect 405660 5370 405688 197678
rect 406580 197674 406608 200086
rect 406476 197668 406528 197674
rect 406476 197610 406528 197616
rect 406568 197668 406620 197674
rect 406568 197610 406620 197616
rect 406384 197532 406436 197538
rect 406384 197474 406436 197480
rect 405648 5364 405700 5370
rect 405648 5306 405700 5312
rect 406016 5228 406068 5234
rect 406016 5170 406068 5176
rect 404820 3528 404872 3534
rect 404820 3470 404872 3476
rect 404832 480 404860 3470
rect 406028 480 406056 5170
rect 406396 3874 406424 197474
rect 406488 14754 406516 197610
rect 406476 14748 406528 14754
rect 406476 14690 406528 14696
rect 407040 5302 407068 200790
rect 407500 197538 407528 200790
rect 407868 197606 407896 200790
rect 407764 197600 407816 197606
rect 407764 197542 407816 197548
rect 407856 197600 407908 197606
rect 407856 197542 407908 197548
rect 407488 197532 407540 197538
rect 407488 197474 407540 197480
rect 407776 17270 407804 197542
rect 408316 197532 408368 197538
rect 408316 197474 408368 197480
rect 407764 17264 407816 17270
rect 407764 17206 407816 17212
rect 408328 8022 408356 197474
rect 408316 8016 408368 8022
rect 408316 7958 408368 7964
rect 407028 5296 407080 5302
rect 407028 5238 407080 5244
rect 408420 5234 408448 200790
rect 408972 197538 409000 200790
rect 409524 197810 409552 200790
rect 409512 197804 409564 197810
rect 409512 197746 409564 197752
rect 409144 197600 409196 197606
rect 409144 197542 409196 197548
rect 408960 197532 409012 197538
rect 408960 197474 409012 197480
rect 408408 5228 408460 5234
rect 408408 5170 408460 5176
rect 407212 5024 407264 5030
rect 407212 4966 407264 4972
rect 406384 3868 406436 3874
rect 406384 3810 406436 3816
rect 407224 480 407252 4966
rect 409156 3806 409184 197542
rect 409696 197532 409748 197538
rect 409696 197474 409748 197480
rect 409708 7954 409736 197474
rect 409696 7948 409748 7954
rect 409696 7890 409748 7896
rect 409800 5166 409828 200790
rect 410444 197538 410472 200790
rect 410904 197606 410932 200790
rect 410892 197600 410944 197606
rect 410892 197542 410944 197548
rect 410432 197532 410484 197538
rect 410432 197474 410484 197480
rect 410984 197532 411036 197538
rect 410984 197474 411036 197480
rect 410996 7886 411024 197474
rect 410984 7880 411036 7886
rect 410984 7822 411036 7828
rect 409604 5160 409656 5166
rect 409604 5102 409656 5108
rect 409788 5160 409840 5166
rect 409788 5102 409840 5108
rect 408408 3800 408460 3806
rect 408408 3742 408460 3748
rect 409144 3800 409196 3806
rect 409144 3742 409196 3748
rect 408420 480 408448 3742
rect 409616 480 409644 5102
rect 410800 5092 410852 5098
rect 410800 5034 410852 5040
rect 410812 480 410840 5034
rect 411088 5030 411116 200926
rect 411746 200790 412128 200818
rect 412298 200790 412588 200818
rect 412758 200790 413048 200818
rect 413310 200790 413784 200818
rect 413862 200790 413968 200818
rect 414322 200790 414704 200818
rect 414874 200790 415164 200818
rect 411168 197600 411220 197606
rect 411168 197542 411220 197548
rect 411076 5024 411128 5030
rect 411076 4966 411128 4972
rect 411180 3738 411208 197542
rect 412100 197538 412128 200790
rect 412560 197742 412588 200790
rect 412548 197736 412600 197742
rect 412548 197678 412600 197684
rect 412088 197532 412140 197538
rect 412088 197474 412140 197480
rect 412548 197532 412600 197538
rect 412548 197474 412600 197480
rect 412560 7818 412588 197474
rect 413020 197402 413048 200790
rect 413008 197396 413060 197402
rect 413008 197338 413060 197344
rect 412548 7812 412600 7818
rect 412548 7754 412600 7760
rect 413756 7750 413784 200790
rect 413836 197396 413888 197402
rect 413836 197338 413888 197344
rect 413744 7744 413796 7750
rect 413744 7686 413796 7692
rect 413848 4962 413876 197338
rect 413100 4956 413152 4962
rect 413100 4898 413152 4904
rect 413836 4956 413888 4962
rect 413836 4898 413888 4904
rect 411168 3732 411220 3738
rect 411168 3674 411220 3680
rect 411904 3460 411956 3466
rect 411904 3402 411956 3408
rect 411916 480 411944 3402
rect 413112 480 413140 4898
rect 413940 3466 413968 200790
rect 414572 198620 414624 198626
rect 414572 198562 414624 198568
rect 414584 190454 414612 198562
rect 414676 197402 414704 200790
rect 415136 200114 415164 200790
rect 415228 200410 415256 200926
rect 415886 200790 416176 200818
rect 416438 200790 416636 200818
rect 416898 200790 417280 200818
rect 417450 200790 417832 200818
rect 417910 200790 418016 200818
rect 418462 200790 418752 200818
rect 419014 200790 419304 200818
rect 415228 200382 415348 200410
rect 415136 200086 415256 200114
rect 414664 197396 414716 197402
rect 414664 197338 414716 197344
rect 414584 190426 414704 190454
rect 414296 4208 414348 4214
rect 414296 4150 414348 4156
rect 413928 3460 413980 3466
rect 413928 3402 413980 3408
rect 414308 480 414336 4150
rect 414676 3534 414704 190426
rect 415228 7682 415256 200086
rect 415320 197674 415348 200382
rect 415308 197668 415360 197674
rect 415308 197610 415360 197616
rect 416148 197402 416176 200790
rect 415308 197396 415360 197402
rect 415308 197338 415360 197344
rect 416136 197396 416188 197402
rect 416136 197338 416188 197344
rect 415216 7676 415268 7682
rect 415216 7618 415268 7624
rect 415320 5098 415348 197338
rect 416608 7614 416636 200790
rect 417252 197470 417280 200790
rect 417240 197464 417292 197470
rect 417240 197406 417292 197412
rect 417804 197402 417832 200790
rect 416688 197396 416740 197402
rect 416688 197338 416740 197344
rect 417424 197396 417476 197402
rect 417424 197338 417476 197344
rect 417792 197396 417844 197402
rect 417792 197338 417844 197344
rect 416596 7608 416648 7614
rect 416596 7550 416648 7556
rect 416700 6914 416728 197338
rect 417436 15978 417464 197338
rect 417424 15972 417476 15978
rect 417424 15914 417476 15920
rect 416608 6886 416728 6914
rect 415308 5092 415360 5098
rect 415308 5034 415360 5040
rect 416608 4962 416636 6886
rect 417988 6186 418016 200790
rect 418724 197402 418752 200790
rect 418896 197532 418948 197538
rect 418896 197474 418948 197480
rect 418804 197464 418856 197470
rect 418804 197406 418856 197412
rect 418068 197396 418120 197402
rect 418068 197338 418120 197344
rect 418712 197396 418764 197402
rect 418712 197338 418764 197344
rect 417976 6180 418028 6186
rect 417976 6122 418028 6128
rect 416596 4956 416648 4962
rect 416596 4898 416648 4904
rect 416688 4888 416740 4894
rect 416688 4830 416740 4836
rect 414664 3528 414716 3534
rect 414664 3470 414716 3476
rect 415492 3528 415544 3534
rect 415492 3470 415544 3476
rect 415504 480 415532 3470
rect 416700 480 416728 4830
rect 418080 4826 418108 197338
rect 418816 6914 418844 197406
rect 418908 14686 418936 197474
rect 419276 190454 419304 200790
rect 419368 198626 419396 200926
rect 420026 200790 420408 200818
rect 419356 198620 419408 198626
rect 419356 198562 419408 198568
rect 420380 198558 420408 200790
rect 420368 198552 420420 198558
rect 420368 198494 420420 198500
rect 420828 198552 420880 198558
rect 420828 198494 420880 198500
rect 419276 190426 419488 190454
rect 418896 14680 418948 14686
rect 418896 14622 418948 14628
rect 418816 6886 419304 6914
rect 417884 4820 417936 4826
rect 417884 4762 417936 4768
rect 418068 4820 418120 4826
rect 418068 4762 418120 4768
rect 417896 480 417924 4762
rect 419276 3602 419304 6886
rect 418988 3596 419040 3602
rect 418988 3538 419040 3544
rect 419264 3596 419316 3602
rect 419264 3538 419316 3544
rect 419000 480 419028 3538
rect 419460 3466 419488 190426
rect 420184 9376 420236 9382
rect 420184 9318 420236 9324
rect 419448 3460 419500 3466
rect 419448 3402 419500 3408
rect 420196 480 420224 9318
rect 420840 3534 420868 198494
rect 421576 20670 421604 506495
rect 421668 46918 421696 508642
rect 421760 86970 421788 508710
rect 421852 126954 421880 508778
rect 421944 458182 421972 509118
rect 422944 508972 422996 508978
rect 422944 508914 422996 508920
rect 421932 458176 421984 458182
rect 421932 458118 421984 458124
rect 422956 206990 422984 508914
rect 422944 206984 422996 206990
rect 422944 206926 422996 206932
rect 422300 197532 422352 197538
rect 422300 197474 422352 197480
rect 421840 126948 421892 126954
rect 421840 126890 421892 126896
rect 421748 86964 421800 86970
rect 421748 86906 421800 86912
rect 421656 46912 421708 46918
rect 421656 46854 421708 46860
rect 421564 20664 421616 20670
rect 421564 20606 421616 20612
rect 422312 16574 422340 197474
rect 424336 73166 424364 510342
rect 425888 509108 425940 509114
rect 425888 509050 425940 509056
rect 424508 509040 424560 509046
rect 424508 508982 424560 508988
rect 424416 508904 424468 508910
rect 424416 508846 424468 508852
rect 424428 167006 424456 508846
rect 424520 245614 424548 508982
rect 425796 507272 425848 507278
rect 425796 507214 425848 507220
rect 425702 506696 425758 506705
rect 425702 506631 425758 506640
rect 424508 245608 424560 245614
rect 424508 245550 424560 245556
rect 424416 167000 424468 167006
rect 424416 166942 424468 166948
rect 424324 73160 424376 73166
rect 424324 73102 424376 73108
rect 425716 60722 425744 506631
rect 425808 113150 425836 507214
rect 425900 299470 425928 509050
rect 426072 507816 426124 507822
rect 426072 507758 426124 507764
rect 425980 507748 426032 507754
rect 425980 507690 426032 507696
rect 425992 405686 426020 507690
rect 426084 485790 426112 507758
rect 429936 507680 429988 507686
rect 429936 507622 429988 507628
rect 428740 507544 428792 507550
rect 428740 507486 428792 507492
rect 428648 507476 428700 507482
rect 428648 507418 428700 507424
rect 428556 507340 428608 507346
rect 428556 507282 428608 507288
rect 428464 507204 428516 507210
rect 428464 507146 428516 507152
rect 426072 485784 426124 485790
rect 426072 485726 426124 485732
rect 425980 405680 426032 405686
rect 425980 405622 426032 405628
rect 425888 299464 425940 299470
rect 425888 299406 425940 299412
rect 425796 113144 425848 113150
rect 425796 113086 425848 113092
rect 428476 100706 428504 507146
rect 428568 153202 428596 507282
rect 428660 193186 428688 507418
rect 428752 233238 428780 507486
rect 429844 507408 429896 507414
rect 429844 507350 429896 507356
rect 428740 233232 428792 233238
rect 428740 233174 428792 233180
rect 429200 198484 429252 198490
rect 429200 198426 429252 198432
rect 428648 193180 428700 193186
rect 428648 193122 428700 193128
rect 428556 153196 428608 153202
rect 428556 153138 428608 153144
rect 428464 100700 428516 100706
rect 428464 100642 428516 100648
rect 425704 60716 425756 60722
rect 425704 60658 425756 60664
rect 423680 19984 423732 19990
rect 423680 19926 423732 19932
rect 423692 16574 423720 19926
rect 422312 16546 422616 16574
rect 423692 16546 423812 16574
rect 421380 7064 421432 7070
rect 421380 7006 421432 7012
rect 420828 3528 420880 3534
rect 420828 3470 420880 3476
rect 421392 480 421420 7006
rect 422588 480 422616 16546
rect 423784 480 423812 16546
rect 427268 9308 427320 9314
rect 427268 9250 427320 9256
rect 424968 7132 425020 7138
rect 424968 7074 425020 7080
rect 424980 480 425008 7074
rect 426164 2984 426216 2990
rect 426164 2926 426216 2932
rect 426176 480 426204 2926
rect 427280 480 427308 9250
rect 428464 7200 428516 7206
rect 428464 7142 428516 7148
rect 428476 480 428504 7142
rect 429212 490 429240 198426
rect 429856 139398 429884 507350
rect 429948 259418 429976 507622
rect 430028 507612 430080 507618
rect 430028 507554 430080 507560
rect 430040 273222 430068 507554
rect 430132 431934 430160 510410
rect 430120 431928 430172 431934
rect 430120 431870 430172 431876
rect 431236 419490 431264 510478
rect 431328 471986 431356 510546
rect 478144 510332 478196 510338
rect 478144 510274 478196 510280
rect 447782 507920 447838 507929
rect 447782 507855 447838 507864
rect 431316 471980 431368 471986
rect 431316 471922 431368 471928
rect 431224 419484 431276 419490
rect 431224 419426 431276 419432
rect 430028 273216 430080 273222
rect 430028 273158 430080 273164
rect 429936 259412 429988 259418
rect 429936 259354 429988 259360
rect 436100 198416 436152 198422
rect 436100 198358 436152 198364
rect 429844 139392 429896 139398
rect 429844 139334 429896 139340
rect 430580 17332 430632 17338
rect 430580 17274 430632 17280
rect 430592 16574 430620 17274
rect 436112 16574 436140 198358
rect 443000 198348 443052 198354
rect 443000 198290 443052 198296
rect 438860 35216 438912 35222
rect 438860 35158 438912 35164
rect 438872 16574 438900 35158
rect 443012 16574 443040 198290
rect 430592 16546 430896 16574
rect 436112 16546 436784 16574
rect 438872 16546 439176 16574
rect 443012 16546 443408 16574
rect 429488 598 429700 626
rect 429488 490 429516 598
rect 371670 -960 371782 480
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376454 -960 376566 480
rect 377650 -960 377762 480
rect 378846 -960 378958 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384734 -960 384846 480
rect 385930 -960 386042 480
rect 387126 -960 387238 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396510 -960 396622 480
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404790 -960 404902 480
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409574 -960 409686 480
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 413070 -960 413182 480
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417854 -960 417966 480
rect 418958 -960 419070 480
rect 420154 -960 420266 480
rect 421350 -960 421462 480
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 426134 -960 426246 480
rect 427238 -960 427350 480
rect 428434 -960 428546 480
rect 429212 462 429516 490
rect 429672 480 429700 598
rect 430868 480 430896 16546
rect 433984 10464 434036 10470
rect 433984 10406 434036 10412
rect 432052 7268 432104 7274
rect 432052 7210 432104 7216
rect 432064 480 432092 7210
rect 433248 3052 433300 3058
rect 433248 2994 433300 3000
rect 433260 480 433288 2994
rect 433996 490 434024 10406
rect 435548 7336 435600 7342
rect 435548 7278 435600 7284
rect 434272 598 434484 626
rect 434272 490 434300 598
rect 429630 -960 429742 480
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 433996 462 434300 490
rect 434456 480 434484 598
rect 435560 480 435588 7278
rect 436756 480 436784 16546
rect 437480 14816 437532 14822
rect 437480 14758 437532 14764
rect 437492 490 437520 14758
rect 437768 598 437980 626
rect 437768 490 437796 598
rect 434414 -960 434526 480
rect 435518 -960 435630 480
rect 436714 -960 436826 480
rect 437492 462 437796 490
rect 437952 480 437980 598
rect 439148 480 439176 16546
rect 442632 16176 442684 16182
rect 442632 16118 442684 16124
rect 441528 13116 441580 13122
rect 441528 13058 441580 13064
rect 440332 3188 440384 3194
rect 440332 3130 440384 3136
rect 440344 480 440372 3130
rect 441540 480 441568 13058
rect 442644 480 442672 16118
rect 443380 490 443408 16546
rect 445760 16108 445812 16114
rect 445760 16050 445812 16056
rect 445024 9172 445076 9178
rect 445024 9114 445076 9120
rect 443656 598 443868 626
rect 443656 490 443684 598
rect 437910 -960 438022 480
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443380 462 443684 490
rect 443840 480 443868 598
rect 445036 480 445064 9114
rect 445772 490 445800 16050
rect 447796 6866 447824 507855
rect 478156 325650 478184 510274
rect 496084 510264 496136 510270
rect 496084 510206 496136 510212
rect 496096 365702 496124 510206
rect 562324 509788 562376 509794
rect 562324 509730 562376 509736
rect 508504 508632 508556 508638
rect 508504 508574 508556 508580
rect 496084 365696 496136 365702
rect 496084 365638 496136 365644
rect 478144 325644 478196 325650
rect 478144 325586 478196 325592
rect 471244 198688 471296 198694
rect 471244 198630 471296 198636
rect 449900 198280 449952 198286
rect 449900 198222 449952 198228
rect 448520 86488 448572 86494
rect 448520 86430 448572 86436
rect 447784 6860 447836 6866
rect 447784 6802 447836 6808
rect 448532 3398 448560 86430
rect 448612 86420 448664 86426
rect 448612 86362 448664 86368
rect 447416 3392 447468 3398
rect 447416 3334 447468 3340
rect 448520 3392 448572 3398
rect 448520 3334 448572 3340
rect 446048 598 446260 626
rect 446048 490 446076 598
rect 443798 -960 443910 480
rect 444994 -960 445106 480
rect 445772 462 446076 490
rect 446232 480 446260 598
rect 447428 480 447456 3334
rect 448624 480 448652 86362
rect 449912 16574 449940 198222
rect 456800 198144 456852 198150
rect 456800 198086 456852 198092
rect 452660 84924 452712 84930
rect 452660 84866 452712 84872
rect 452672 16574 452700 84866
rect 449912 16546 450952 16574
rect 452672 16546 453344 16574
rect 449808 3392 449860 3398
rect 449808 3334 449860 3340
rect 449820 480 449848 3334
rect 450924 480 450952 16546
rect 452108 5636 452160 5642
rect 452108 5578 452160 5584
rect 452120 480 452148 5578
rect 453316 480 453344 16546
rect 455696 5704 455748 5710
rect 455696 5646 455748 5652
rect 454500 3256 454552 3262
rect 454500 3198 454552 3204
rect 454512 480 454540 3198
rect 455708 480 455736 5646
rect 456812 3398 456840 198086
rect 467840 198076 467892 198082
rect 467840 198018 467892 198024
rect 467104 197940 467156 197946
rect 467104 197882 467156 197888
rect 456892 87644 456944 87650
rect 456892 87586 456944 87592
rect 456800 3392 456852 3398
rect 456800 3334 456852 3340
rect 456904 480 456932 87586
rect 463700 25560 463752 25566
rect 463700 25502 463752 25508
rect 463712 16574 463740 25502
rect 467116 16574 467144 197882
rect 467852 16574 467880 198018
rect 470600 44872 470652 44878
rect 470600 44814 470652 44820
rect 463712 16546 464016 16574
rect 467116 16546 467236 16574
rect 467852 16546 468248 16574
rect 460388 9240 460440 9246
rect 460388 9182 460440 9188
rect 459192 5772 459244 5778
rect 459192 5714 459244 5720
rect 458088 3392 458140 3398
rect 458088 3334 458140 3340
rect 458100 480 458128 3334
rect 459204 480 459232 5714
rect 460400 480 460428 9182
rect 462780 5840 462832 5846
rect 462780 5782 462832 5788
rect 461584 3324 461636 3330
rect 461584 3266 461636 3272
rect 461596 480 461624 3266
rect 462792 480 462820 5782
rect 463988 480 464016 16546
rect 467104 16244 467156 16250
rect 467104 16186 467156 16192
rect 466276 5908 466328 5914
rect 466276 5850 466328 5856
rect 465172 3120 465224 3126
rect 465172 3062 465224 3068
rect 465184 480 465212 3062
rect 466288 480 466316 5850
rect 467116 2802 467144 16186
rect 467208 2990 467236 16546
rect 467196 2984 467248 2990
rect 467196 2926 467248 2932
rect 467116 2774 467512 2802
rect 467484 480 467512 2774
rect 468220 490 468248 16546
rect 469864 5976 469916 5982
rect 469864 5918 469916 5924
rect 468496 598 468708 626
rect 468496 490 468524 598
rect 446190 -960 446302 480
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 452078 -960 452190 480
rect 453274 -960 453386 480
rect 454470 -960 454582 480
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 460358 -960 460470 480
rect 461554 -960 461666 480
rect 462750 -960 462862 480
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 466246 -960 466358 480
rect 467442 -960 467554 480
rect 468220 462 468524 490
rect 468680 480 468708 598
rect 469876 480 469904 5918
rect 470612 490 470640 44814
rect 471256 3058 471284 198630
rect 490564 198620 490616 198626
rect 490564 198562 490616 198568
rect 482376 198212 482428 198218
rect 482376 198154 482428 198160
rect 474740 198008 474792 198014
rect 474740 197950 474792 197956
rect 472624 197872 472676 197878
rect 472624 197814 472676 197820
rect 472256 4140 472308 4146
rect 472256 4082 472308 4088
rect 471244 3052 471296 3058
rect 471244 2994 471296 3000
rect 470888 598 471100 626
rect 470888 490 470916 598
rect 468638 -960 468750 480
rect 469834 -960 469946 480
rect 470612 462 470916 490
rect 471072 480 471100 598
rect 472268 480 472296 4082
rect 472636 3126 472664 197814
rect 474004 197600 474056 197606
rect 474004 197542 474056 197548
rect 473912 10328 473964 10334
rect 473912 10270 473964 10276
rect 473452 6112 473504 6118
rect 473452 6054 473504 6060
rect 472624 3120 472676 3126
rect 472624 3062 472676 3068
rect 473464 480 473492 6054
rect 473924 626 473952 10270
rect 474016 3194 474044 197542
rect 474752 16574 474780 197950
rect 478144 197804 478196 197810
rect 478144 197746 478196 197752
rect 478156 16574 478184 197746
rect 479524 197736 479576 197742
rect 479524 197678 479576 197684
rect 474752 16546 475792 16574
rect 478156 16546 478276 16574
rect 474004 3188 474056 3194
rect 474004 3130 474056 3136
rect 473924 598 474136 626
rect 474108 490 474136 598
rect 474384 598 474596 626
rect 474384 490 474412 598
rect 471030 -960 471142 480
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 474108 462 474412 490
rect 474568 480 474596 598
rect 475764 480 475792 16546
rect 478052 9104 478104 9110
rect 478052 9046 478104 9052
rect 476948 6044 477000 6050
rect 476948 5986 477000 5992
rect 476960 480 476988 5986
rect 478064 3482 478092 9046
rect 478064 3454 478184 3482
rect 478156 480 478184 3454
rect 478248 3262 478276 16546
rect 479340 4072 479392 4078
rect 479340 4014 479392 4020
rect 478236 3256 478288 3262
rect 478236 3198 478288 3204
rect 479352 480 479380 4014
rect 479536 3330 479564 197678
rect 482284 197532 482336 197538
rect 482284 197474 482336 197480
rect 482100 10396 482152 10402
rect 482100 10338 482152 10344
rect 480536 9036 480588 9042
rect 480536 8978 480588 8984
rect 479524 3324 479576 3330
rect 479524 3266 479576 3272
rect 480548 480 480576 8978
rect 481732 6792 481784 6798
rect 481732 6734 481784 6740
rect 481744 480 481772 6734
rect 482112 626 482140 10338
rect 482296 6914 482324 197474
rect 482388 9042 482416 198154
rect 486424 197396 486476 197402
rect 486424 197338 486476 197344
rect 485780 86352 485832 86358
rect 485780 86294 485832 86300
rect 485792 16574 485820 86294
rect 485792 16546 486372 16574
rect 484032 16040 484084 16046
rect 484032 15982 484084 15988
rect 482376 9036 482428 9042
rect 482376 8978 482428 8984
rect 482204 6886 482324 6914
rect 482204 3398 482232 6886
rect 482192 3392 482244 3398
rect 482192 3334 482244 3340
rect 482112 598 482416 626
rect 482388 490 482416 598
rect 482664 598 482876 626
rect 482664 490 482692 598
rect 474526 -960 474638 480
rect 475722 -960 475834 480
rect 476918 -960 477030 480
rect 478114 -960 478226 480
rect 479310 -960 479422 480
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482388 462 482692 490
rect 482848 480 482876 598
rect 484044 480 484072 15982
rect 485228 6724 485280 6730
rect 485228 6666 485280 6672
rect 485240 480 485268 6666
rect 486344 3482 486372 16546
rect 486436 4078 486464 197338
rect 489920 196784 489972 196790
rect 489920 196726 489972 196732
rect 487160 11824 487212 11830
rect 487160 11766 487212 11772
rect 486424 4072 486476 4078
rect 486424 4014 486476 4020
rect 486344 3454 486464 3482
rect 486436 480 486464 3454
rect 487172 490 487200 11766
rect 488816 6656 488868 6662
rect 488816 6598 488868 6604
rect 487448 598 487660 626
rect 487448 490 487476 598
rect 482806 -960 482918 480
rect 484002 -960 484114 480
rect 485198 -960 485310 480
rect 486394 -960 486506 480
rect 487172 462 487476 490
rect 487632 480 487660 598
rect 488828 480 488856 6598
rect 489932 4146 489960 196726
rect 490576 16574 490604 198562
rect 505100 196716 505152 196722
rect 505100 196658 505152 196664
rect 500960 89004 501012 89010
rect 500960 88946 501012 88952
rect 499580 26920 499632 26926
rect 499580 26862 499632 26868
rect 492680 21412 492732 21418
rect 492680 21354 492732 21360
rect 492692 16574 492720 21354
rect 496820 17264 496872 17270
rect 496820 17206 496872 17212
rect 496832 16574 496860 17206
rect 499592 16574 499620 26862
rect 500972 16574 501000 88946
rect 503720 84856 503772 84862
rect 503720 84798 503772 84804
rect 490576 16546 490788 16574
rect 492692 16546 493088 16574
rect 496832 16546 497136 16574
rect 499592 16546 500632 16574
rect 500972 16546 501368 16574
rect 490012 14748 490064 14754
rect 490012 14690 490064 14696
rect 489920 4140 489972 4146
rect 489920 4082 489972 4088
rect 490024 3482 490052 14690
rect 490760 4214 490788 16546
rect 492312 6588 492364 6594
rect 492312 6530 492364 6536
rect 490748 4208 490800 4214
rect 490748 4150 490800 4156
rect 491116 4140 491168 4146
rect 491116 4082 491168 4088
rect 489932 3454 490052 3482
rect 489932 480 489960 3454
rect 491128 480 491156 4082
rect 492324 480 492352 6530
rect 493060 490 493088 16546
rect 494704 11756 494756 11762
rect 494704 11698 494756 11704
rect 493336 598 493548 626
rect 493336 490 493364 598
rect 487590 -960 487702 480
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 491086 -960 491198 480
rect 492282 -960 492394 480
rect 493060 462 493364 490
rect 493520 480 493548 598
rect 494716 480 494744 11698
rect 495900 6520 495952 6526
rect 495900 6462 495952 6468
rect 495912 480 495940 6462
rect 497108 480 497136 16546
rect 498200 8968 498252 8974
rect 498200 8910 498252 8916
rect 498212 480 498240 8910
rect 499396 6452 499448 6458
rect 499396 6394 499448 6400
rect 499408 480 499436 6394
rect 500604 480 500632 16546
rect 501340 490 501368 16546
rect 502984 6384 503036 6390
rect 502984 6326 503036 6332
rect 501616 598 501828 626
rect 501616 490 501644 598
rect 493478 -960 493590 480
rect 494674 -960 494786 480
rect 495870 -960 495982 480
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 499366 -960 499478 480
rect 500562 -960 500674 480
rect 501340 462 501644 490
rect 501800 480 501828 598
rect 502996 480 503024 6326
rect 503732 490 503760 84798
rect 505112 16574 505140 196658
rect 506480 86284 506532 86290
rect 506480 86226 506532 86232
rect 506492 16574 506520 86226
rect 508516 33114 508544 508574
rect 562336 379506 562364 509730
rect 573364 508428 573416 508434
rect 573364 508370 573416 508376
rect 562324 379500 562376 379506
rect 562324 379442 562376 379448
rect 573376 353258 573404 508370
rect 580264 507136 580316 507142
rect 580264 507078 580316 507084
rect 580172 485784 580224 485790
rect 580172 485726 580224 485732
rect 580184 484673 580212 485726
rect 580170 484664 580226 484673
rect 580170 484599 580226 484608
rect 580172 471980 580224 471986
rect 580172 471922 580224 471928
rect 580184 471481 580212 471922
rect 580170 471472 580226 471481
rect 580170 471407 580226 471416
rect 580172 458176 580224 458182
rect 580170 458144 580172 458153
rect 580224 458144 580226 458153
rect 580170 458079 580226 458088
rect 580172 431928 580224 431934
rect 580172 431870 580224 431876
rect 580184 431633 580212 431870
rect 580170 431624 580226 431633
rect 580170 431559 580226 431568
rect 579712 419484 579764 419490
rect 579712 419426 579764 419432
rect 579724 418305 579752 419426
rect 579710 418296 579766 418305
rect 579710 418231 579766 418240
rect 579804 405680 579856 405686
rect 579804 405622 579856 405628
rect 579816 404977 579844 405622
rect 579802 404968 579858 404977
rect 579802 404903 579858 404912
rect 579804 379500 579856 379506
rect 579804 379442 579856 379448
rect 579816 378457 579844 379442
rect 579802 378448 579858 378457
rect 579802 378383 579858 378392
rect 580172 365696 580224 365702
rect 580172 365638 580224 365644
rect 580184 365129 580212 365638
rect 580170 365120 580226 365129
rect 580170 365055 580226 365064
rect 573364 353252 573416 353258
rect 573364 353194 573416 353200
rect 579620 353252 579672 353258
rect 579620 353194 579672 353200
rect 579632 351937 579660 353194
rect 579618 351928 579674 351937
rect 579618 351863 579674 351872
rect 580172 325644 580224 325650
rect 580172 325586 580224 325592
rect 580184 325281 580212 325586
rect 580170 325272 580226 325281
rect 580170 325207 580226 325216
rect 580172 299464 580224 299470
rect 580172 299406 580224 299412
rect 580184 298761 580212 299406
rect 580170 298752 580226 298761
rect 580170 298687 580226 298696
rect 580172 273216 580224 273222
rect 580172 273158 580224 273164
rect 580184 272241 580212 273158
rect 580170 272232 580226 272241
rect 580170 272167 580226 272176
rect 579620 259412 579672 259418
rect 579620 259354 579672 259360
rect 579632 258913 579660 259354
rect 579618 258904 579674 258913
rect 579618 258839 579674 258848
rect 580172 245608 580224 245614
rect 580170 245576 580172 245585
rect 580224 245576 580226 245585
rect 580170 245511 580226 245520
rect 580172 233232 580224 233238
rect 580172 233174 580224 233180
rect 580184 232393 580212 233174
rect 580170 232384 580226 232393
rect 580170 232319 580226 232328
rect 580172 206984 580224 206990
rect 580172 206926 580224 206932
rect 580184 205737 580212 206926
rect 580170 205728 580226 205737
rect 580170 205663 580226 205672
rect 516140 196648 516192 196654
rect 516140 196590 516192 196596
rect 508504 33108 508556 33114
rect 508504 33050 508556 33056
rect 514760 24132 514812 24138
rect 514760 24074 514812 24080
rect 505112 16546 505416 16574
rect 506492 16546 507256 16574
rect 504008 598 504220 626
rect 504008 490 504036 598
rect 501758 -960 501870 480
rect 502954 -960 503066 480
rect 503732 462 504036 490
rect 504192 480 504220 598
rect 505388 480 505416 16546
rect 506480 6316 506532 6322
rect 506480 6258 506532 6264
rect 506492 480 506520 6258
rect 507228 490 507256 16546
rect 508872 15904 508924 15910
rect 508872 15846 508924 15852
rect 507504 598 507716 626
rect 507504 490 507532 598
rect 504150 -960 504262 480
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 507228 462 507532 490
rect 507688 480 507716 598
rect 508884 480 508912 15846
rect 511264 14680 511316 14686
rect 511264 14622 511316 14628
rect 510068 6248 510120 6254
rect 510068 6190 510120 6196
rect 510080 480 510108 6190
rect 511276 480 511304 14622
rect 513564 14612 513616 14618
rect 513564 14554 513616 14560
rect 512460 4276 512512 4282
rect 512460 4218 512512 4224
rect 512472 480 512500 4218
rect 513576 480 513604 14554
rect 514772 480 514800 24074
rect 516152 16574 516180 196590
rect 580172 193180 580224 193186
rect 580172 193122 580224 193128
rect 580184 192545 580212 193122
rect 580170 192536 580226 192545
rect 580170 192471 580226 192480
rect 580276 179217 580304 507078
rect 580448 506728 580500 506734
rect 580448 506670 580500 506676
rect 580356 506660 580408 506666
rect 580356 506602 580408 506608
rect 580368 219065 580396 506602
rect 580460 312089 580488 506670
rect 580446 312080 580502 312089
rect 580446 312015 580502 312024
rect 580354 219056 580410 219065
rect 580354 218991 580410 219000
rect 580262 179208 580318 179217
rect 580262 179143 580318 179152
rect 580172 167000 580224 167006
rect 580172 166942 580224 166948
rect 580184 165889 580212 166942
rect 580170 165880 580226 165889
rect 580170 165815 580226 165824
rect 580172 153196 580224 153202
rect 580172 153138 580224 153144
rect 580184 152697 580212 153138
rect 580170 152688 580226 152697
rect 580170 152623 580226 152632
rect 580172 139392 580224 139398
rect 580170 139360 580172 139369
rect 580224 139360 580226 139369
rect 580170 139295 580226 139304
rect 580172 126948 580224 126954
rect 580172 126890 580224 126896
rect 580184 126041 580212 126890
rect 580170 126032 580226 126041
rect 580170 125967 580226 125976
rect 579804 113144 579856 113150
rect 579804 113086 579856 113092
rect 579816 112849 579844 113086
rect 579802 112840 579858 112849
rect 579802 112775 579858 112784
rect 580172 100700 580224 100706
rect 580172 100642 580224 100648
rect 580184 99521 580212 100642
rect 580170 99512 580226 99521
rect 580170 99447 580226 99456
rect 580172 86964 580224 86970
rect 580172 86906 580224 86912
rect 580184 86193 580212 86906
rect 580170 86184 580226 86193
rect 580170 86119 580226 86128
rect 580172 73160 580224 73166
rect 580172 73102 580224 73108
rect 580184 73001 580212 73102
rect 580170 72992 580226 73001
rect 580170 72927 580226 72936
rect 580172 60716 580224 60722
rect 580172 60658 580224 60664
rect 580184 59673 580212 60658
rect 580170 59664 580226 59673
rect 580170 59599 580226 59608
rect 580172 46912 580224 46918
rect 580172 46854 580224 46860
rect 580184 46345 580212 46854
rect 580170 46336 580226 46345
rect 580170 46271 580226 46280
rect 580170 33144 580226 33153
rect 580170 33079 580172 33088
rect 580224 33079 580226 33088
rect 580172 33050 580224 33056
rect 521660 22772 521712 22778
rect 521660 22714 521712 22720
rect 521672 16574 521700 22714
rect 579988 20664 580040 20670
rect 579988 20606 580040 20612
rect 580000 19825 580028 20606
rect 579986 19816 580042 19825
rect 579986 19751 580042 19760
rect 516152 16546 517192 16574
rect 521672 16546 521884 16574
rect 515956 4344 516008 4350
rect 515956 4286 516008 4292
rect 515968 480 515996 4286
rect 517164 480 517192 16546
rect 520280 14476 520332 14482
rect 520280 14418 520332 14424
rect 518348 9036 518400 9042
rect 518348 8978 518400 8984
rect 518360 480 518388 8978
rect 519544 4412 519596 4418
rect 519544 4354 519596 4360
rect 519556 480 519584 4354
rect 520292 490 520320 14418
rect 520568 598 520780 626
rect 520568 490 520596 598
rect 507646 -960 507758 480
rect 508842 -960 508954 480
rect 510038 -960 510150 480
rect 511234 -960 511346 480
rect 512430 -960 512542 480
rect 513534 -960 513646 480
rect 514730 -960 514842 480
rect 515926 -960 516038 480
rect 517122 -960 517234 480
rect 518318 -960 518430 480
rect 519514 -960 519626 480
rect 520292 462 520596 490
rect 520752 480 520780 598
rect 521856 480 521884 16546
rect 525432 15972 525484 15978
rect 525432 15914 525484 15920
rect 522304 14544 522356 14550
rect 522304 14486 522356 14492
rect 522316 2990 522344 14486
rect 523040 4480 523092 4486
rect 523040 4422 523092 4428
rect 522304 2984 522356 2990
rect 522304 2926 522356 2932
rect 523052 480 523080 4422
rect 524236 2984 524288 2990
rect 524236 2926 524288 2932
rect 524248 480 524276 2926
rect 525444 480 525472 15914
rect 538404 8288 538456 8294
rect 538404 8230 538456 8236
rect 534908 7540 534960 7546
rect 534908 7482 534960 7488
rect 531320 7472 531372 7478
rect 531320 7414 531372 7420
rect 527824 7404 527876 7410
rect 527824 7346 527876 7352
rect 526628 4548 526680 4554
rect 526628 4490 526680 4496
rect 526640 480 526668 4490
rect 527836 480 527864 7346
rect 530124 4616 530176 4622
rect 530124 4558 530176 4564
rect 529020 2916 529072 2922
rect 529020 2858 529072 2864
rect 529032 480 529060 2858
rect 530136 480 530164 4558
rect 531332 480 531360 7414
rect 533712 4684 533764 4690
rect 533712 4626 533764 4632
rect 532516 4004 532568 4010
rect 532516 3946 532568 3952
rect 532528 480 532556 3946
rect 533724 480 533752 4626
rect 534920 480 534948 7482
rect 537208 4752 537260 4758
rect 537208 4694 537260 4700
rect 536104 3052 536156 3058
rect 536104 2994 536156 3000
rect 536116 480 536144 2994
rect 537220 480 537248 4694
rect 538416 480 538444 8230
rect 541992 8220 542044 8226
rect 541992 8162 542044 8168
rect 540796 5500 540848 5506
rect 540796 5442 540848 5448
rect 539600 3936 539652 3942
rect 539600 3878 539652 3884
rect 539612 480 539640 3878
rect 540808 480 540836 5442
rect 542004 480 542032 8162
rect 545488 8152 545540 8158
rect 545488 8094 545540 8100
rect 544384 5432 544436 5438
rect 544384 5374 544436 5380
rect 543188 3120 543240 3126
rect 543188 3062 543240 3068
rect 543200 480 543228 3062
rect 544396 480 544424 5374
rect 545500 480 545528 8094
rect 549076 8084 549128 8090
rect 549076 8026 549128 8032
rect 547880 5364 547932 5370
rect 547880 5306 547932 5312
rect 546684 3868 546736 3874
rect 546684 3810 546736 3816
rect 546696 480 546724 3810
rect 547892 480 547920 5306
rect 549088 480 549116 8026
rect 552664 8016 552716 8022
rect 552664 7958 552716 7964
rect 551468 5296 551520 5302
rect 551468 5238 551520 5244
rect 550272 3188 550324 3194
rect 550272 3130 550324 3136
rect 550284 480 550312 3130
rect 551480 480 551508 5238
rect 552676 480 552704 7958
rect 556160 7948 556212 7954
rect 556160 7890 556212 7896
rect 554964 5228 555016 5234
rect 554964 5170 555016 5176
rect 553768 3800 553820 3806
rect 553768 3742 553820 3748
rect 553780 480 553808 3742
rect 554976 480 555004 5170
rect 556172 480 556200 7890
rect 559748 7880 559800 7886
rect 559748 7822 559800 7828
rect 558552 5160 558604 5166
rect 558552 5102 558604 5108
rect 557356 3256 557408 3262
rect 557356 3198 557408 3204
rect 557368 480 557396 3198
rect 558564 480 558592 5102
rect 559760 480 559788 7822
rect 563244 7812 563296 7818
rect 563244 7754 563296 7760
rect 562048 5024 562100 5030
rect 562048 4966 562100 4972
rect 560852 3732 560904 3738
rect 560852 3674 560904 3680
rect 560864 480 560892 3674
rect 562060 480 562088 4966
rect 563256 480 563284 7754
rect 566832 7744 566884 7750
rect 566832 7686 566884 7692
rect 565636 5092 565688 5098
rect 565636 5034 565688 5040
rect 564440 3324 564492 3330
rect 564440 3266 564492 3272
rect 564452 480 564480 3266
rect 565648 480 565676 5034
rect 566844 480 566872 7686
rect 570328 7676 570380 7682
rect 570328 7618 570380 7624
rect 569132 4956 569184 4962
rect 569132 4898 569184 4904
rect 568028 3664 568080 3670
rect 568028 3606 568080 3612
rect 568040 480 568068 3606
rect 569144 480 569172 4898
rect 570340 480 570368 7618
rect 573916 7608 573968 7614
rect 573916 7550 573968 7556
rect 572720 4888 572772 4894
rect 572720 4830 572772 4836
rect 571524 3392 571576 3398
rect 571524 3334 571576 3340
rect 571536 480 571564 3334
rect 572732 480 572760 4830
rect 573928 480 573956 7550
rect 580172 6860 580224 6866
rect 580172 6802 580224 6808
rect 580184 6633 580212 6802
rect 580170 6624 580226 6633
rect 580170 6559 580226 6568
rect 577412 6180 577464 6186
rect 577412 6122 577464 6128
rect 576308 4820 576360 4826
rect 576308 4762 576360 4768
rect 575112 3596 575164 3602
rect 575112 3538 575164 3544
rect 575124 480 575152 3538
rect 576320 480 576348 4762
rect 577424 480 577452 6122
rect 582196 4140 582248 4146
rect 582196 4082 582248 4088
rect 578608 4072 578660 4078
rect 578608 4014 578660 4020
rect 578620 480 578648 4014
rect 581000 3460 581052 3466
rect 581000 3402 581052 3408
rect 581012 480 581040 3402
rect 582208 480 582236 4082
rect 583392 3528 583444 3534
rect 583392 3470 583444 3476
rect 583404 480 583432 3470
rect 520710 -960 520822 480
rect 521814 -960 521926 480
rect 523010 -960 523122 480
rect 524206 -960 524318 480
rect 525402 -960 525514 480
rect 526598 -960 526710 480
rect 527794 -960 527906 480
rect 528990 -960 529102 480
rect 530094 -960 530206 480
rect 531290 -960 531402 480
rect 532486 -960 532598 480
rect 533682 -960 533794 480
rect 534878 -960 534990 480
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538374 -960 538486 480
rect 539570 -960 539682 480
rect 540766 -960 540878 480
rect 541962 -960 542074 480
rect 543158 -960 543270 480
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546654 -960 546766 480
rect 547850 -960 547962 480
rect 549046 -960 549158 480
rect 550242 -960 550354 480
rect 551438 -960 551550 480
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554934 -960 555046 480
rect 556130 -960 556242 480
rect 557326 -960 557438 480
rect 558522 -960 558634 480
rect 559718 -960 559830 480
rect 560822 -960 560934 480
rect 562018 -960 562130 480
rect 563214 -960 563326 480
rect 564410 -960 564522 480
rect 565606 -960 565718 480
rect 566802 -960 566914 480
rect 567998 -960 568110 480
rect 569102 -960 569214 480
rect 570298 -960 570410 480
rect 571494 -960 571606 480
rect 572690 -960 572802 480
rect 573886 -960 573998 480
rect 575082 -960 575194 480
rect 576278 -960 576390 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 3422 684256 3478 684312
rect 3514 671200 3570 671256
rect 3422 658144 3478 658200
rect 3422 632068 3424 632088
rect 3424 632068 3476 632088
rect 3476 632068 3478 632088
rect 3422 632032 3478 632068
rect 3146 619112 3202 619168
rect 3238 606056 3294 606112
rect 3330 579944 3386 580000
rect 3422 566888 3478 566944
rect 3422 553832 3478 553888
rect 3422 527856 3478 527912
rect 3422 514820 3478 514856
rect 3422 514800 3424 514820
rect 3424 514800 3476 514820
rect 3476 514800 3478 514820
rect 3422 509224 3478 509280
rect 3146 501744 3202 501800
rect 3330 475668 3332 475688
rect 3332 475668 3384 475688
rect 3384 475668 3386 475688
rect 3330 475632 3386 475668
rect 2778 462576 2834 462632
rect 3330 449520 3386 449576
rect 3330 423580 3332 423600
rect 3332 423580 3384 423600
rect 3384 423580 3386 423600
rect 3330 423544 3386 423580
rect 2778 410488 2834 410544
rect 3330 397432 3386 397488
rect 3054 371320 3110 371376
rect 2778 358436 2780 358456
rect 2780 358436 2832 358456
rect 2832 358436 2834 358456
rect 2778 358400 2834 358436
rect 3330 345344 3386 345400
rect 3330 319232 3386 319288
rect 3330 306176 3386 306232
rect 2870 293120 2926 293176
rect 3238 267144 3294 267200
rect 3330 254088 3386 254144
rect 3330 214956 3332 214976
rect 3332 214956 3384 214976
rect 3384 214956 3386 214976
rect 3330 214920 3386 214956
rect 3054 201864 3110 201920
rect 2778 188844 2780 188864
rect 2780 188844 2832 188864
rect 2832 188844 2834 188864
rect 2778 188808 2834 188844
rect 3330 162832 3386 162888
rect 3054 58520 3110 58576
rect 2870 32408 2926 32464
rect 3606 241032 3662 241088
rect 3606 149776 3662 149832
rect 3514 136720 3570 136776
rect 3514 110608 3570 110664
rect 3514 97552 3570 97608
rect 3514 84632 3570 84688
rect 3514 71612 3516 71632
rect 3516 71612 3568 71632
rect 3568 71612 3570 71632
rect 3514 71576 3570 71612
rect 3514 45500 3516 45520
rect 3516 45500 3568 45520
rect 3568 45500 3570 45520
rect 3514 45464 3570 45500
rect 3514 19352 3570 19408
rect 3422 6432 3478 6488
rect 166814 507864 166870 507920
rect 580170 697176 580226 697232
rect 580170 683848 580226 683904
rect 580170 670656 580226 670712
rect 580170 644000 580226 644056
rect 580170 630808 580226 630864
rect 580170 617480 580226 617536
rect 579802 590960 579858 591016
rect 580170 577632 580226 577688
rect 579802 564304 579858 564360
rect 580170 537784 580226 537840
rect 580170 524476 580226 524512
rect 580170 524456 580172 524476
rect 580172 524456 580224 524476
rect 580224 524456 580226 524476
rect 580170 511264 580226 511320
rect 416962 509224 417018 509280
rect 171598 507320 171654 507376
rect 178406 507320 178462 507376
rect 421562 506504 421618 506560
rect 425702 506640 425758 506696
rect 447782 507864 447838 507920
rect 580170 484608 580226 484664
rect 580170 471416 580226 471472
rect 580170 458124 580172 458144
rect 580172 458124 580224 458144
rect 580224 458124 580226 458144
rect 580170 458088 580226 458124
rect 580170 431568 580226 431624
rect 579710 418240 579766 418296
rect 579802 404912 579858 404968
rect 579802 378392 579858 378448
rect 580170 365064 580226 365120
rect 579618 351872 579674 351928
rect 580170 325216 580226 325272
rect 580170 298696 580226 298752
rect 580170 272176 580226 272232
rect 579618 258848 579674 258904
rect 580170 245556 580172 245576
rect 580172 245556 580224 245576
rect 580224 245556 580226 245576
rect 580170 245520 580226 245556
rect 580170 232328 580226 232384
rect 580170 205672 580226 205728
rect 580170 192480 580226 192536
rect 580446 312024 580502 312080
rect 580354 219000 580410 219056
rect 580262 179152 580318 179208
rect 580170 165824 580226 165880
rect 580170 152632 580226 152688
rect 580170 139340 580172 139360
rect 580172 139340 580224 139360
rect 580224 139340 580226 139360
rect 580170 139304 580226 139340
rect 580170 125976 580226 126032
rect 579802 112784 579858 112840
rect 580170 99456 580226 99512
rect 580170 86128 580226 86184
rect 580170 72936 580226 72992
rect 580170 59608 580226 59664
rect 580170 46280 580226 46336
rect 580170 33108 580226 33144
rect 580170 33088 580172 33108
rect 580172 33088 580224 33108
rect 580224 33088 580226 33108
rect 579986 19760 580042 19816
rect 580170 6568 580226 6624
<< metal3 >>
rect -960 697220 480 697460
rect 580165 697234 580231 697237
rect 583520 697234 584960 697324
rect 580165 697232 584960 697234
rect 580165 697176 580170 697232
rect 580226 697176 584960 697232
rect 580165 697174 584960 697176
rect 580165 697171 580231 697174
rect 583520 697084 584960 697174
rect -960 684314 480 684404
rect 3417 684314 3483 684317
rect -960 684312 3483 684314
rect -960 684256 3422 684312
rect 3478 684256 3483 684312
rect -960 684254 3483 684256
rect -960 684164 480 684254
rect 3417 684251 3483 684254
rect 580165 683906 580231 683909
rect 583520 683906 584960 683996
rect 580165 683904 584960 683906
rect 580165 683848 580170 683904
rect 580226 683848 584960 683904
rect 580165 683846 584960 683848
rect 580165 683843 580231 683846
rect 583520 683756 584960 683846
rect -960 671258 480 671348
rect 3509 671258 3575 671261
rect -960 671256 3575 671258
rect -960 671200 3514 671256
rect 3570 671200 3575 671256
rect -960 671198 3575 671200
rect -960 671108 480 671198
rect 3509 671195 3575 671198
rect 580165 670714 580231 670717
rect 583520 670714 584960 670804
rect 580165 670712 584960 670714
rect 580165 670656 580170 670712
rect 580226 670656 584960 670712
rect 580165 670654 584960 670656
rect 580165 670651 580231 670654
rect 583520 670564 584960 670654
rect -960 658202 480 658292
rect 3417 658202 3483 658205
rect -960 658200 3483 658202
rect -960 658144 3422 658200
rect 3478 658144 3483 658200
rect -960 658142 3483 658144
rect -960 658052 480 658142
rect 3417 658139 3483 658142
rect 583520 657236 584960 657476
rect -960 644996 480 645236
rect 580165 644058 580231 644061
rect 583520 644058 584960 644148
rect 580165 644056 584960 644058
rect 580165 644000 580170 644056
rect 580226 644000 584960 644056
rect 580165 643998 584960 644000
rect 580165 643995 580231 643998
rect 583520 643908 584960 643998
rect -960 632090 480 632180
rect 3417 632090 3483 632093
rect -960 632088 3483 632090
rect -960 632032 3422 632088
rect 3478 632032 3483 632088
rect -960 632030 3483 632032
rect -960 631940 480 632030
rect 3417 632027 3483 632030
rect 580165 630866 580231 630869
rect 583520 630866 584960 630956
rect 580165 630864 584960 630866
rect 580165 630808 580170 630864
rect 580226 630808 584960 630864
rect 580165 630806 584960 630808
rect 580165 630803 580231 630806
rect 583520 630716 584960 630806
rect -960 619170 480 619260
rect 3141 619170 3207 619173
rect -960 619168 3207 619170
rect -960 619112 3146 619168
rect 3202 619112 3207 619168
rect -960 619110 3207 619112
rect -960 619020 480 619110
rect 3141 619107 3207 619110
rect 580165 617538 580231 617541
rect 583520 617538 584960 617628
rect 580165 617536 584960 617538
rect 580165 617480 580170 617536
rect 580226 617480 584960 617536
rect 580165 617478 584960 617480
rect 580165 617475 580231 617478
rect 583520 617388 584960 617478
rect -960 606114 480 606204
rect 3233 606114 3299 606117
rect -960 606112 3299 606114
rect -960 606056 3238 606112
rect 3294 606056 3299 606112
rect -960 606054 3299 606056
rect -960 605964 480 606054
rect 3233 606051 3299 606054
rect 583520 604060 584960 604300
rect -960 592908 480 593148
rect 579797 591018 579863 591021
rect 583520 591018 584960 591108
rect 579797 591016 584960 591018
rect 579797 590960 579802 591016
rect 579858 590960 584960 591016
rect 579797 590958 584960 590960
rect 579797 590955 579863 590958
rect 583520 590868 584960 590958
rect -960 580002 480 580092
rect 3325 580002 3391 580005
rect -960 580000 3391 580002
rect -960 579944 3330 580000
rect 3386 579944 3391 580000
rect -960 579942 3391 579944
rect -960 579852 480 579942
rect 3325 579939 3391 579942
rect 580165 577690 580231 577693
rect 583520 577690 584960 577780
rect 580165 577688 584960 577690
rect 580165 577632 580170 577688
rect 580226 577632 584960 577688
rect 580165 577630 584960 577632
rect 580165 577627 580231 577630
rect 583520 577540 584960 577630
rect -960 566946 480 567036
rect 3417 566946 3483 566949
rect -960 566944 3483 566946
rect -960 566888 3422 566944
rect 3478 566888 3483 566944
rect -960 566886 3483 566888
rect -960 566796 480 566886
rect 3417 566883 3483 566886
rect 579797 564362 579863 564365
rect 583520 564362 584960 564452
rect 579797 564360 584960 564362
rect 579797 564304 579802 564360
rect 579858 564304 584960 564360
rect 579797 564302 584960 564304
rect 579797 564299 579863 564302
rect 583520 564212 584960 564302
rect -960 553890 480 553980
rect 3417 553890 3483 553893
rect -960 553888 3483 553890
rect -960 553832 3422 553888
rect 3478 553832 3483 553888
rect -960 553830 3483 553832
rect -960 553740 480 553830
rect 3417 553827 3483 553830
rect 583520 551020 584960 551260
rect -960 540684 480 540924
rect 580165 537842 580231 537845
rect 583520 537842 584960 537932
rect 580165 537840 584960 537842
rect 580165 537784 580170 537840
rect 580226 537784 584960 537840
rect 580165 537782 584960 537784
rect 580165 537779 580231 537782
rect 583520 537692 584960 537782
rect -960 527914 480 528004
rect 3417 527914 3483 527917
rect -960 527912 3483 527914
rect -960 527856 3422 527912
rect 3478 527856 3483 527912
rect -960 527854 3483 527856
rect -960 527764 480 527854
rect 3417 527851 3483 527854
rect 580165 524514 580231 524517
rect 583520 524514 584960 524604
rect 580165 524512 584960 524514
rect 580165 524456 580170 524512
rect 580226 524456 584960 524512
rect 580165 524454 584960 524456
rect 580165 524451 580231 524454
rect 583520 524364 584960 524454
rect -960 514858 480 514948
rect 3417 514858 3483 514861
rect -960 514856 3483 514858
rect -960 514800 3422 514856
rect 3478 514800 3483 514856
rect -960 514798 3483 514800
rect -960 514708 480 514798
rect 3417 514795 3483 514798
rect 580165 511322 580231 511325
rect 583520 511322 584960 511412
rect 580165 511320 584960 511322
rect 580165 511264 580170 511320
rect 580226 511264 584960 511320
rect 580165 511262 584960 511264
rect 580165 511259 580231 511262
rect 583520 511172 584960 511262
rect 3417 509282 3483 509285
rect 416957 509282 417023 509285
rect 3417 509280 417023 509282
rect 3417 509224 3422 509280
rect 3478 509224 416962 509280
rect 417018 509224 417023 509280
rect 3417 509222 417023 509224
rect 3417 509219 3483 509222
rect 416957 509219 417023 509222
rect 166809 507922 166875 507925
rect 447777 507922 447843 507925
rect 166809 507920 447843 507922
rect 166809 507864 166814 507920
rect 166870 507864 447782 507920
rect 447838 507864 447843 507920
rect 166809 507862 447843 507864
rect 166809 507859 166875 507862
rect 447777 507859 447843 507862
rect 171593 507378 171659 507381
rect 178401 507378 178467 507381
rect 171593 507376 176026 507378
rect 171593 507320 171598 507376
rect 171654 507320 176026 507376
rect 171593 507318 176026 507320
rect 171593 507315 171659 507318
rect 175966 506562 176026 507318
rect 178401 507376 180810 507378
rect 178401 507320 178406 507376
rect 178462 507320 180810 507376
rect 178401 507318 180810 507320
rect 178401 507315 178467 507318
rect 180750 506698 180810 507318
rect 425697 506698 425763 506701
rect 180750 506696 425763 506698
rect 180750 506640 425702 506696
rect 425758 506640 425763 506696
rect 180750 506638 425763 506640
rect 425697 506635 425763 506638
rect 421557 506562 421623 506565
rect 175966 506560 421623 506562
rect 175966 506504 421562 506560
rect 421618 506504 421623 506560
rect 175966 506502 421623 506504
rect 421557 506499 421623 506502
rect -960 501802 480 501892
rect 3141 501802 3207 501805
rect -960 501800 3207 501802
rect -960 501744 3146 501800
rect 3202 501744 3207 501800
rect -960 501742 3207 501744
rect -960 501652 480 501742
rect 3141 501739 3207 501742
rect 583520 497844 584960 498084
rect -960 488596 480 488836
rect 580165 484666 580231 484669
rect 583520 484666 584960 484756
rect 580165 484664 584960 484666
rect 580165 484608 580170 484664
rect 580226 484608 584960 484664
rect 580165 484606 584960 484608
rect 580165 484603 580231 484606
rect 583520 484516 584960 484606
rect -960 475690 480 475780
rect 3325 475690 3391 475693
rect -960 475688 3391 475690
rect -960 475632 3330 475688
rect 3386 475632 3391 475688
rect -960 475630 3391 475632
rect -960 475540 480 475630
rect 3325 475627 3391 475630
rect 580165 471474 580231 471477
rect 583520 471474 584960 471564
rect 580165 471472 584960 471474
rect 580165 471416 580170 471472
rect 580226 471416 584960 471472
rect 580165 471414 584960 471416
rect 580165 471411 580231 471414
rect 583520 471324 584960 471414
rect -960 462634 480 462724
rect 2773 462634 2839 462637
rect -960 462632 2839 462634
rect -960 462576 2778 462632
rect 2834 462576 2839 462632
rect -960 462574 2839 462576
rect -960 462484 480 462574
rect 2773 462571 2839 462574
rect 580165 458146 580231 458149
rect 583520 458146 584960 458236
rect 580165 458144 584960 458146
rect 580165 458088 580170 458144
rect 580226 458088 584960 458144
rect 580165 458086 584960 458088
rect 580165 458083 580231 458086
rect 583520 457996 584960 458086
rect -960 449578 480 449668
rect 3325 449578 3391 449581
rect -960 449576 3391 449578
rect -960 449520 3330 449576
rect 3386 449520 3391 449576
rect -960 449518 3391 449520
rect -960 449428 480 449518
rect 3325 449515 3391 449518
rect 583520 444668 584960 444908
rect -960 436508 480 436748
rect 580165 431626 580231 431629
rect 583520 431626 584960 431716
rect 580165 431624 584960 431626
rect 580165 431568 580170 431624
rect 580226 431568 584960 431624
rect 580165 431566 584960 431568
rect 580165 431563 580231 431566
rect 583520 431476 584960 431566
rect -960 423602 480 423692
rect 3325 423602 3391 423605
rect -960 423600 3391 423602
rect -960 423544 3330 423600
rect 3386 423544 3391 423600
rect -960 423542 3391 423544
rect -960 423452 480 423542
rect 3325 423539 3391 423542
rect 579705 418298 579771 418301
rect 583520 418298 584960 418388
rect 579705 418296 584960 418298
rect 579705 418240 579710 418296
rect 579766 418240 584960 418296
rect 579705 418238 584960 418240
rect 579705 418235 579771 418238
rect 583520 418148 584960 418238
rect -960 410546 480 410636
rect 2773 410546 2839 410549
rect -960 410544 2839 410546
rect -960 410488 2778 410544
rect 2834 410488 2839 410544
rect -960 410486 2839 410488
rect -960 410396 480 410486
rect 2773 410483 2839 410486
rect 579797 404970 579863 404973
rect 583520 404970 584960 405060
rect 579797 404968 584960 404970
rect 579797 404912 579802 404968
rect 579858 404912 584960 404968
rect 579797 404910 584960 404912
rect 579797 404907 579863 404910
rect 583520 404820 584960 404910
rect -960 397490 480 397580
rect 3325 397490 3391 397493
rect -960 397488 3391 397490
rect -960 397432 3330 397488
rect 3386 397432 3391 397488
rect -960 397430 3391 397432
rect -960 397340 480 397430
rect 3325 397427 3391 397430
rect 583520 391628 584960 391868
rect -960 384284 480 384524
rect 579797 378450 579863 378453
rect 583520 378450 584960 378540
rect 579797 378448 584960 378450
rect 579797 378392 579802 378448
rect 579858 378392 584960 378448
rect 579797 378390 584960 378392
rect 579797 378387 579863 378390
rect 583520 378300 584960 378390
rect -960 371378 480 371468
rect 3049 371378 3115 371381
rect -960 371376 3115 371378
rect -960 371320 3054 371376
rect 3110 371320 3115 371376
rect -960 371318 3115 371320
rect -960 371228 480 371318
rect 3049 371315 3115 371318
rect 580165 365122 580231 365125
rect 583520 365122 584960 365212
rect 580165 365120 584960 365122
rect 580165 365064 580170 365120
rect 580226 365064 584960 365120
rect 580165 365062 584960 365064
rect 580165 365059 580231 365062
rect 583520 364972 584960 365062
rect -960 358458 480 358548
rect 2773 358458 2839 358461
rect -960 358456 2839 358458
rect -960 358400 2778 358456
rect 2834 358400 2839 358456
rect -960 358398 2839 358400
rect -960 358308 480 358398
rect 2773 358395 2839 358398
rect 579613 351930 579679 351933
rect 583520 351930 584960 352020
rect 579613 351928 584960 351930
rect 579613 351872 579618 351928
rect 579674 351872 584960 351928
rect 579613 351870 584960 351872
rect 579613 351867 579679 351870
rect 583520 351780 584960 351870
rect -960 345402 480 345492
rect 3325 345402 3391 345405
rect -960 345400 3391 345402
rect -960 345344 3330 345400
rect 3386 345344 3391 345400
rect -960 345342 3391 345344
rect -960 345252 480 345342
rect 3325 345339 3391 345342
rect 583520 338452 584960 338692
rect -960 332196 480 332436
rect 580165 325274 580231 325277
rect 583520 325274 584960 325364
rect 580165 325272 584960 325274
rect 580165 325216 580170 325272
rect 580226 325216 584960 325272
rect 580165 325214 584960 325216
rect 580165 325211 580231 325214
rect 583520 325124 584960 325214
rect -960 319290 480 319380
rect 3325 319290 3391 319293
rect -960 319288 3391 319290
rect -960 319232 3330 319288
rect 3386 319232 3391 319288
rect -960 319230 3391 319232
rect -960 319140 480 319230
rect 3325 319227 3391 319230
rect 580441 312082 580507 312085
rect 583520 312082 584960 312172
rect 580441 312080 584960 312082
rect 580441 312024 580446 312080
rect 580502 312024 584960 312080
rect 580441 312022 584960 312024
rect 580441 312019 580507 312022
rect 583520 311932 584960 312022
rect -960 306234 480 306324
rect 3325 306234 3391 306237
rect -960 306232 3391 306234
rect -960 306176 3330 306232
rect 3386 306176 3391 306232
rect -960 306174 3391 306176
rect -960 306084 480 306174
rect 3325 306171 3391 306174
rect 580165 298754 580231 298757
rect 583520 298754 584960 298844
rect 580165 298752 584960 298754
rect 580165 298696 580170 298752
rect 580226 298696 584960 298752
rect 580165 298694 584960 298696
rect 580165 298691 580231 298694
rect 583520 298604 584960 298694
rect -960 293178 480 293268
rect 2865 293178 2931 293181
rect -960 293176 2931 293178
rect -960 293120 2870 293176
rect 2926 293120 2931 293176
rect -960 293118 2931 293120
rect -960 293028 480 293118
rect 2865 293115 2931 293118
rect 583520 285276 584960 285516
rect -960 279972 480 280212
rect 580165 272234 580231 272237
rect 583520 272234 584960 272324
rect 580165 272232 584960 272234
rect 580165 272176 580170 272232
rect 580226 272176 584960 272232
rect 580165 272174 584960 272176
rect 580165 272171 580231 272174
rect 583520 272084 584960 272174
rect -960 267202 480 267292
rect 3233 267202 3299 267205
rect -960 267200 3299 267202
rect -960 267144 3238 267200
rect 3294 267144 3299 267200
rect -960 267142 3299 267144
rect -960 267052 480 267142
rect 3233 267139 3299 267142
rect 579613 258906 579679 258909
rect 583520 258906 584960 258996
rect 579613 258904 584960 258906
rect 579613 258848 579618 258904
rect 579674 258848 584960 258904
rect 579613 258846 584960 258848
rect 579613 258843 579679 258846
rect 583520 258756 584960 258846
rect -960 254146 480 254236
rect 3325 254146 3391 254149
rect -960 254144 3391 254146
rect -960 254088 3330 254144
rect 3386 254088 3391 254144
rect -960 254086 3391 254088
rect -960 253996 480 254086
rect 3325 254083 3391 254086
rect 580165 245578 580231 245581
rect 583520 245578 584960 245668
rect 580165 245576 584960 245578
rect 580165 245520 580170 245576
rect 580226 245520 584960 245576
rect 580165 245518 584960 245520
rect 580165 245515 580231 245518
rect 583520 245428 584960 245518
rect -960 241090 480 241180
rect 3601 241090 3667 241093
rect -960 241088 3667 241090
rect -960 241032 3606 241088
rect 3662 241032 3667 241088
rect -960 241030 3667 241032
rect -960 240940 480 241030
rect 3601 241027 3667 241030
rect 580165 232386 580231 232389
rect 583520 232386 584960 232476
rect 580165 232384 584960 232386
rect 580165 232328 580170 232384
rect 580226 232328 584960 232384
rect 580165 232326 584960 232328
rect 580165 232323 580231 232326
rect 583520 232236 584960 232326
rect -960 227884 480 228124
rect 580349 219058 580415 219061
rect 583520 219058 584960 219148
rect 580349 219056 584960 219058
rect 580349 219000 580354 219056
rect 580410 219000 584960 219056
rect 580349 218998 584960 219000
rect 580349 218995 580415 218998
rect 583520 218908 584960 218998
rect -960 214978 480 215068
rect 3325 214978 3391 214981
rect -960 214976 3391 214978
rect -960 214920 3330 214976
rect 3386 214920 3391 214976
rect -960 214918 3391 214920
rect -960 214828 480 214918
rect 3325 214915 3391 214918
rect 580165 205730 580231 205733
rect 583520 205730 584960 205820
rect 580165 205728 584960 205730
rect 580165 205672 580170 205728
rect 580226 205672 584960 205728
rect 580165 205670 584960 205672
rect 580165 205667 580231 205670
rect 583520 205580 584960 205670
rect -960 201922 480 202012
rect 3049 201922 3115 201925
rect -960 201920 3115 201922
rect -960 201864 3054 201920
rect 3110 201864 3115 201920
rect -960 201862 3115 201864
rect -960 201772 480 201862
rect 3049 201859 3115 201862
rect 580165 192538 580231 192541
rect 583520 192538 584960 192628
rect 580165 192536 584960 192538
rect 580165 192480 580170 192536
rect 580226 192480 584960 192536
rect 580165 192478 584960 192480
rect 580165 192475 580231 192478
rect 583520 192388 584960 192478
rect -960 188866 480 188956
rect 2773 188866 2839 188869
rect -960 188864 2839 188866
rect -960 188808 2778 188864
rect 2834 188808 2839 188864
rect -960 188806 2839 188808
rect -960 188716 480 188806
rect 2773 188803 2839 188806
rect 580257 179210 580323 179213
rect 583520 179210 584960 179300
rect 580257 179208 584960 179210
rect 580257 179152 580262 179208
rect 580318 179152 584960 179208
rect 580257 179150 584960 179152
rect 580257 179147 580323 179150
rect 583520 179060 584960 179150
rect -960 175796 480 176036
rect 580165 165882 580231 165885
rect 583520 165882 584960 165972
rect 580165 165880 584960 165882
rect 580165 165824 580170 165880
rect 580226 165824 584960 165880
rect 580165 165822 584960 165824
rect 580165 165819 580231 165822
rect 583520 165732 584960 165822
rect -960 162890 480 162980
rect 3325 162890 3391 162893
rect -960 162888 3391 162890
rect -960 162832 3330 162888
rect 3386 162832 3391 162888
rect -960 162830 3391 162832
rect -960 162740 480 162830
rect 3325 162827 3391 162830
rect 580165 152690 580231 152693
rect 583520 152690 584960 152780
rect 580165 152688 584960 152690
rect 580165 152632 580170 152688
rect 580226 152632 584960 152688
rect 580165 152630 584960 152632
rect 580165 152627 580231 152630
rect 583520 152540 584960 152630
rect -960 149834 480 149924
rect 3601 149834 3667 149837
rect -960 149832 3667 149834
rect -960 149776 3606 149832
rect 3662 149776 3667 149832
rect -960 149774 3667 149776
rect -960 149684 480 149774
rect 3601 149771 3667 149774
rect 580165 139362 580231 139365
rect 583520 139362 584960 139452
rect 580165 139360 584960 139362
rect 580165 139304 580170 139360
rect 580226 139304 584960 139360
rect 580165 139302 584960 139304
rect 580165 139299 580231 139302
rect 583520 139212 584960 139302
rect -960 136778 480 136868
rect 3509 136778 3575 136781
rect -960 136776 3575 136778
rect -960 136720 3514 136776
rect 3570 136720 3575 136776
rect -960 136718 3575 136720
rect -960 136628 480 136718
rect 3509 136715 3575 136718
rect 580165 126034 580231 126037
rect 583520 126034 584960 126124
rect 580165 126032 584960 126034
rect 580165 125976 580170 126032
rect 580226 125976 584960 126032
rect 580165 125974 584960 125976
rect 580165 125971 580231 125974
rect 583520 125884 584960 125974
rect -960 123572 480 123812
rect 579797 112842 579863 112845
rect 583520 112842 584960 112932
rect 579797 112840 584960 112842
rect 579797 112784 579802 112840
rect 579858 112784 584960 112840
rect 579797 112782 584960 112784
rect 579797 112779 579863 112782
rect 583520 112692 584960 112782
rect -960 110666 480 110756
rect 3509 110666 3575 110669
rect -960 110664 3575 110666
rect -960 110608 3514 110664
rect 3570 110608 3575 110664
rect -960 110606 3575 110608
rect -960 110516 480 110606
rect 3509 110603 3575 110606
rect 580165 99514 580231 99517
rect 583520 99514 584960 99604
rect 580165 99512 584960 99514
rect 580165 99456 580170 99512
rect 580226 99456 584960 99512
rect 580165 99454 584960 99456
rect 580165 99451 580231 99454
rect 583520 99364 584960 99454
rect -960 97610 480 97700
rect 3509 97610 3575 97613
rect -960 97608 3575 97610
rect -960 97552 3514 97608
rect 3570 97552 3575 97608
rect -960 97550 3575 97552
rect -960 97460 480 97550
rect 3509 97547 3575 97550
rect 580165 86186 580231 86189
rect 583520 86186 584960 86276
rect 580165 86184 584960 86186
rect 580165 86128 580170 86184
rect 580226 86128 584960 86184
rect 580165 86126 584960 86128
rect 580165 86123 580231 86126
rect 583520 86036 584960 86126
rect -960 84690 480 84780
rect 3509 84690 3575 84693
rect -960 84688 3575 84690
rect -960 84632 3514 84688
rect 3570 84632 3575 84688
rect -960 84630 3575 84632
rect -960 84540 480 84630
rect 3509 84627 3575 84630
rect 580165 72994 580231 72997
rect 583520 72994 584960 73084
rect 580165 72992 584960 72994
rect 580165 72936 580170 72992
rect 580226 72936 584960 72992
rect 580165 72934 584960 72936
rect 580165 72931 580231 72934
rect 583520 72844 584960 72934
rect -960 71634 480 71724
rect 3509 71634 3575 71637
rect -960 71632 3575 71634
rect -960 71576 3514 71632
rect 3570 71576 3575 71632
rect -960 71574 3575 71576
rect -960 71484 480 71574
rect 3509 71571 3575 71574
rect 580165 59666 580231 59669
rect 583520 59666 584960 59756
rect 580165 59664 584960 59666
rect 580165 59608 580170 59664
rect 580226 59608 584960 59664
rect 580165 59606 584960 59608
rect 580165 59603 580231 59606
rect 583520 59516 584960 59606
rect -960 58578 480 58668
rect 3049 58578 3115 58581
rect -960 58576 3115 58578
rect -960 58520 3054 58576
rect 3110 58520 3115 58576
rect -960 58518 3115 58520
rect -960 58428 480 58518
rect 3049 58515 3115 58518
rect 580165 46338 580231 46341
rect 583520 46338 584960 46428
rect 580165 46336 584960 46338
rect 580165 46280 580170 46336
rect 580226 46280 584960 46336
rect 580165 46278 584960 46280
rect 580165 46275 580231 46278
rect 583520 46188 584960 46278
rect -960 45522 480 45612
rect 3509 45522 3575 45525
rect -960 45520 3575 45522
rect -960 45464 3514 45520
rect 3570 45464 3575 45520
rect -960 45462 3575 45464
rect -960 45372 480 45462
rect 3509 45459 3575 45462
rect 580165 33146 580231 33149
rect 583520 33146 584960 33236
rect 580165 33144 584960 33146
rect 580165 33088 580170 33144
rect 580226 33088 584960 33144
rect 580165 33086 584960 33088
rect 580165 33083 580231 33086
rect 583520 32996 584960 33086
rect -960 32466 480 32556
rect 2865 32466 2931 32469
rect -960 32464 2931 32466
rect -960 32408 2870 32464
rect 2926 32408 2931 32464
rect -960 32406 2931 32408
rect -960 32316 480 32406
rect 2865 32403 2931 32406
rect 579981 19818 580047 19821
rect 583520 19818 584960 19908
rect 579981 19816 584960 19818
rect 579981 19760 579986 19816
rect 580042 19760 584960 19816
rect 579981 19758 584960 19760
rect 579981 19755 580047 19758
rect 583520 19668 584960 19758
rect -960 19410 480 19500
rect 3509 19410 3575 19413
rect -960 19408 3575 19410
rect -960 19352 3514 19408
rect 3570 19352 3575 19408
rect -960 19350 3575 19352
rect -960 19260 480 19350
rect 3509 19347 3575 19350
rect 580165 6626 580231 6629
rect 583520 6626 584960 6716
rect 580165 6624 584960 6626
rect -960 6490 480 6580
rect 580165 6568 580170 6624
rect 580226 6568 584960 6624
rect 580165 6566 584960 6568
rect 580165 6563 580231 6566
rect 3417 6490 3483 6493
rect -960 6488 3483 6490
rect -960 6432 3422 6488
rect 3478 6432 3483 6488
rect 583520 6476 584960 6566
rect -960 6430 3483 6432
rect -960 6340 480 6430
rect 3417 6427 3483 6430
<< metal4 >>
rect -8726 711558 -8106 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 -8106 711558
rect -8726 711238 -8106 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 -8106 711238
rect -8726 680614 -8106 711002
rect -8726 680378 -8694 680614
rect -8458 680378 -8374 680614
rect -8138 680378 -8106 680614
rect -8726 680294 -8106 680378
rect -8726 680058 -8694 680294
rect -8458 680058 -8374 680294
rect -8138 680058 -8106 680294
rect -8726 644614 -8106 680058
rect -8726 644378 -8694 644614
rect -8458 644378 -8374 644614
rect -8138 644378 -8106 644614
rect -8726 644294 -8106 644378
rect -8726 644058 -8694 644294
rect -8458 644058 -8374 644294
rect -8138 644058 -8106 644294
rect -8726 608614 -8106 644058
rect -8726 608378 -8694 608614
rect -8458 608378 -8374 608614
rect -8138 608378 -8106 608614
rect -8726 608294 -8106 608378
rect -8726 608058 -8694 608294
rect -8458 608058 -8374 608294
rect -8138 608058 -8106 608294
rect -8726 572614 -8106 608058
rect -8726 572378 -8694 572614
rect -8458 572378 -8374 572614
rect -8138 572378 -8106 572614
rect -8726 572294 -8106 572378
rect -8726 572058 -8694 572294
rect -8458 572058 -8374 572294
rect -8138 572058 -8106 572294
rect -8726 536614 -8106 572058
rect -8726 536378 -8694 536614
rect -8458 536378 -8374 536614
rect -8138 536378 -8106 536614
rect -8726 536294 -8106 536378
rect -8726 536058 -8694 536294
rect -8458 536058 -8374 536294
rect -8138 536058 -8106 536294
rect -8726 500614 -8106 536058
rect -8726 500378 -8694 500614
rect -8458 500378 -8374 500614
rect -8138 500378 -8106 500614
rect -8726 500294 -8106 500378
rect -8726 500058 -8694 500294
rect -8458 500058 -8374 500294
rect -8138 500058 -8106 500294
rect -8726 464614 -8106 500058
rect -8726 464378 -8694 464614
rect -8458 464378 -8374 464614
rect -8138 464378 -8106 464614
rect -8726 464294 -8106 464378
rect -8726 464058 -8694 464294
rect -8458 464058 -8374 464294
rect -8138 464058 -8106 464294
rect -8726 428614 -8106 464058
rect -8726 428378 -8694 428614
rect -8458 428378 -8374 428614
rect -8138 428378 -8106 428614
rect -8726 428294 -8106 428378
rect -8726 428058 -8694 428294
rect -8458 428058 -8374 428294
rect -8138 428058 -8106 428294
rect -8726 392614 -8106 428058
rect -8726 392378 -8694 392614
rect -8458 392378 -8374 392614
rect -8138 392378 -8106 392614
rect -8726 392294 -8106 392378
rect -8726 392058 -8694 392294
rect -8458 392058 -8374 392294
rect -8138 392058 -8106 392294
rect -8726 356614 -8106 392058
rect -8726 356378 -8694 356614
rect -8458 356378 -8374 356614
rect -8138 356378 -8106 356614
rect -8726 356294 -8106 356378
rect -8726 356058 -8694 356294
rect -8458 356058 -8374 356294
rect -8138 356058 -8106 356294
rect -8726 320614 -8106 356058
rect -8726 320378 -8694 320614
rect -8458 320378 -8374 320614
rect -8138 320378 -8106 320614
rect -8726 320294 -8106 320378
rect -8726 320058 -8694 320294
rect -8458 320058 -8374 320294
rect -8138 320058 -8106 320294
rect -8726 284614 -8106 320058
rect -8726 284378 -8694 284614
rect -8458 284378 -8374 284614
rect -8138 284378 -8106 284614
rect -8726 284294 -8106 284378
rect -8726 284058 -8694 284294
rect -8458 284058 -8374 284294
rect -8138 284058 -8106 284294
rect -8726 248614 -8106 284058
rect -8726 248378 -8694 248614
rect -8458 248378 -8374 248614
rect -8138 248378 -8106 248614
rect -8726 248294 -8106 248378
rect -8726 248058 -8694 248294
rect -8458 248058 -8374 248294
rect -8138 248058 -8106 248294
rect -8726 212614 -8106 248058
rect -8726 212378 -8694 212614
rect -8458 212378 -8374 212614
rect -8138 212378 -8106 212614
rect -8726 212294 -8106 212378
rect -8726 212058 -8694 212294
rect -8458 212058 -8374 212294
rect -8138 212058 -8106 212294
rect -8726 176614 -8106 212058
rect -8726 176378 -8694 176614
rect -8458 176378 -8374 176614
rect -8138 176378 -8106 176614
rect -8726 176294 -8106 176378
rect -8726 176058 -8694 176294
rect -8458 176058 -8374 176294
rect -8138 176058 -8106 176294
rect -8726 140614 -8106 176058
rect -8726 140378 -8694 140614
rect -8458 140378 -8374 140614
rect -8138 140378 -8106 140614
rect -8726 140294 -8106 140378
rect -8726 140058 -8694 140294
rect -8458 140058 -8374 140294
rect -8138 140058 -8106 140294
rect -8726 104614 -8106 140058
rect -8726 104378 -8694 104614
rect -8458 104378 -8374 104614
rect -8138 104378 -8106 104614
rect -8726 104294 -8106 104378
rect -8726 104058 -8694 104294
rect -8458 104058 -8374 104294
rect -8138 104058 -8106 104294
rect -8726 68614 -8106 104058
rect -8726 68378 -8694 68614
rect -8458 68378 -8374 68614
rect -8138 68378 -8106 68614
rect -8726 68294 -8106 68378
rect -8726 68058 -8694 68294
rect -8458 68058 -8374 68294
rect -8138 68058 -8106 68294
rect -8726 32614 -8106 68058
rect -8726 32378 -8694 32614
rect -8458 32378 -8374 32614
rect -8138 32378 -8106 32614
rect -8726 32294 -8106 32378
rect -8726 32058 -8694 32294
rect -8458 32058 -8374 32294
rect -8138 32058 -8106 32294
rect -8726 -7066 -8106 32058
rect -7766 710598 -7146 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 -7146 710598
rect -7766 710278 -7146 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 -7146 710278
rect -7766 698614 -7146 710042
rect 12954 710598 13574 711590
rect 12954 710362 12986 710598
rect 13222 710362 13306 710598
rect 13542 710362 13574 710598
rect 12954 710278 13574 710362
rect 12954 710042 12986 710278
rect 13222 710042 13306 710278
rect 13542 710042 13574 710278
rect -7766 698378 -7734 698614
rect -7498 698378 -7414 698614
rect -7178 698378 -7146 698614
rect -7766 698294 -7146 698378
rect -7766 698058 -7734 698294
rect -7498 698058 -7414 698294
rect -7178 698058 -7146 698294
rect -7766 662614 -7146 698058
rect -7766 662378 -7734 662614
rect -7498 662378 -7414 662614
rect -7178 662378 -7146 662614
rect -7766 662294 -7146 662378
rect -7766 662058 -7734 662294
rect -7498 662058 -7414 662294
rect -7178 662058 -7146 662294
rect -7766 626614 -7146 662058
rect -7766 626378 -7734 626614
rect -7498 626378 -7414 626614
rect -7178 626378 -7146 626614
rect -7766 626294 -7146 626378
rect -7766 626058 -7734 626294
rect -7498 626058 -7414 626294
rect -7178 626058 -7146 626294
rect -7766 590614 -7146 626058
rect -7766 590378 -7734 590614
rect -7498 590378 -7414 590614
rect -7178 590378 -7146 590614
rect -7766 590294 -7146 590378
rect -7766 590058 -7734 590294
rect -7498 590058 -7414 590294
rect -7178 590058 -7146 590294
rect -7766 554614 -7146 590058
rect -7766 554378 -7734 554614
rect -7498 554378 -7414 554614
rect -7178 554378 -7146 554614
rect -7766 554294 -7146 554378
rect -7766 554058 -7734 554294
rect -7498 554058 -7414 554294
rect -7178 554058 -7146 554294
rect -7766 518614 -7146 554058
rect -7766 518378 -7734 518614
rect -7498 518378 -7414 518614
rect -7178 518378 -7146 518614
rect -7766 518294 -7146 518378
rect -7766 518058 -7734 518294
rect -7498 518058 -7414 518294
rect -7178 518058 -7146 518294
rect -7766 482614 -7146 518058
rect -7766 482378 -7734 482614
rect -7498 482378 -7414 482614
rect -7178 482378 -7146 482614
rect -7766 482294 -7146 482378
rect -7766 482058 -7734 482294
rect -7498 482058 -7414 482294
rect -7178 482058 -7146 482294
rect -7766 446614 -7146 482058
rect -7766 446378 -7734 446614
rect -7498 446378 -7414 446614
rect -7178 446378 -7146 446614
rect -7766 446294 -7146 446378
rect -7766 446058 -7734 446294
rect -7498 446058 -7414 446294
rect -7178 446058 -7146 446294
rect -7766 410614 -7146 446058
rect -7766 410378 -7734 410614
rect -7498 410378 -7414 410614
rect -7178 410378 -7146 410614
rect -7766 410294 -7146 410378
rect -7766 410058 -7734 410294
rect -7498 410058 -7414 410294
rect -7178 410058 -7146 410294
rect -7766 374614 -7146 410058
rect -7766 374378 -7734 374614
rect -7498 374378 -7414 374614
rect -7178 374378 -7146 374614
rect -7766 374294 -7146 374378
rect -7766 374058 -7734 374294
rect -7498 374058 -7414 374294
rect -7178 374058 -7146 374294
rect -7766 338614 -7146 374058
rect -7766 338378 -7734 338614
rect -7498 338378 -7414 338614
rect -7178 338378 -7146 338614
rect -7766 338294 -7146 338378
rect -7766 338058 -7734 338294
rect -7498 338058 -7414 338294
rect -7178 338058 -7146 338294
rect -7766 302614 -7146 338058
rect -7766 302378 -7734 302614
rect -7498 302378 -7414 302614
rect -7178 302378 -7146 302614
rect -7766 302294 -7146 302378
rect -7766 302058 -7734 302294
rect -7498 302058 -7414 302294
rect -7178 302058 -7146 302294
rect -7766 266614 -7146 302058
rect -7766 266378 -7734 266614
rect -7498 266378 -7414 266614
rect -7178 266378 -7146 266614
rect -7766 266294 -7146 266378
rect -7766 266058 -7734 266294
rect -7498 266058 -7414 266294
rect -7178 266058 -7146 266294
rect -7766 230614 -7146 266058
rect -7766 230378 -7734 230614
rect -7498 230378 -7414 230614
rect -7178 230378 -7146 230614
rect -7766 230294 -7146 230378
rect -7766 230058 -7734 230294
rect -7498 230058 -7414 230294
rect -7178 230058 -7146 230294
rect -7766 194614 -7146 230058
rect -7766 194378 -7734 194614
rect -7498 194378 -7414 194614
rect -7178 194378 -7146 194614
rect -7766 194294 -7146 194378
rect -7766 194058 -7734 194294
rect -7498 194058 -7414 194294
rect -7178 194058 -7146 194294
rect -7766 158614 -7146 194058
rect -7766 158378 -7734 158614
rect -7498 158378 -7414 158614
rect -7178 158378 -7146 158614
rect -7766 158294 -7146 158378
rect -7766 158058 -7734 158294
rect -7498 158058 -7414 158294
rect -7178 158058 -7146 158294
rect -7766 122614 -7146 158058
rect -7766 122378 -7734 122614
rect -7498 122378 -7414 122614
rect -7178 122378 -7146 122614
rect -7766 122294 -7146 122378
rect -7766 122058 -7734 122294
rect -7498 122058 -7414 122294
rect -7178 122058 -7146 122294
rect -7766 86614 -7146 122058
rect -7766 86378 -7734 86614
rect -7498 86378 -7414 86614
rect -7178 86378 -7146 86614
rect -7766 86294 -7146 86378
rect -7766 86058 -7734 86294
rect -7498 86058 -7414 86294
rect -7178 86058 -7146 86294
rect -7766 50614 -7146 86058
rect -7766 50378 -7734 50614
rect -7498 50378 -7414 50614
rect -7178 50378 -7146 50614
rect -7766 50294 -7146 50378
rect -7766 50058 -7734 50294
rect -7498 50058 -7414 50294
rect -7178 50058 -7146 50294
rect -7766 14614 -7146 50058
rect -7766 14378 -7734 14614
rect -7498 14378 -7414 14614
rect -7178 14378 -7146 14614
rect -7766 14294 -7146 14378
rect -7766 14058 -7734 14294
rect -7498 14058 -7414 14294
rect -7178 14058 -7146 14294
rect -7766 -6106 -7146 14058
rect -6806 709638 -6186 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 -6186 709638
rect -6806 709318 -6186 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 -6186 709318
rect -6806 676894 -6186 709082
rect -6806 676658 -6774 676894
rect -6538 676658 -6454 676894
rect -6218 676658 -6186 676894
rect -6806 676574 -6186 676658
rect -6806 676338 -6774 676574
rect -6538 676338 -6454 676574
rect -6218 676338 -6186 676574
rect -6806 640894 -6186 676338
rect -6806 640658 -6774 640894
rect -6538 640658 -6454 640894
rect -6218 640658 -6186 640894
rect -6806 640574 -6186 640658
rect -6806 640338 -6774 640574
rect -6538 640338 -6454 640574
rect -6218 640338 -6186 640574
rect -6806 604894 -6186 640338
rect -6806 604658 -6774 604894
rect -6538 604658 -6454 604894
rect -6218 604658 -6186 604894
rect -6806 604574 -6186 604658
rect -6806 604338 -6774 604574
rect -6538 604338 -6454 604574
rect -6218 604338 -6186 604574
rect -6806 568894 -6186 604338
rect -6806 568658 -6774 568894
rect -6538 568658 -6454 568894
rect -6218 568658 -6186 568894
rect -6806 568574 -6186 568658
rect -6806 568338 -6774 568574
rect -6538 568338 -6454 568574
rect -6218 568338 -6186 568574
rect -6806 532894 -6186 568338
rect -6806 532658 -6774 532894
rect -6538 532658 -6454 532894
rect -6218 532658 -6186 532894
rect -6806 532574 -6186 532658
rect -6806 532338 -6774 532574
rect -6538 532338 -6454 532574
rect -6218 532338 -6186 532574
rect -6806 496894 -6186 532338
rect -6806 496658 -6774 496894
rect -6538 496658 -6454 496894
rect -6218 496658 -6186 496894
rect -6806 496574 -6186 496658
rect -6806 496338 -6774 496574
rect -6538 496338 -6454 496574
rect -6218 496338 -6186 496574
rect -6806 460894 -6186 496338
rect -6806 460658 -6774 460894
rect -6538 460658 -6454 460894
rect -6218 460658 -6186 460894
rect -6806 460574 -6186 460658
rect -6806 460338 -6774 460574
rect -6538 460338 -6454 460574
rect -6218 460338 -6186 460574
rect -6806 424894 -6186 460338
rect -6806 424658 -6774 424894
rect -6538 424658 -6454 424894
rect -6218 424658 -6186 424894
rect -6806 424574 -6186 424658
rect -6806 424338 -6774 424574
rect -6538 424338 -6454 424574
rect -6218 424338 -6186 424574
rect -6806 388894 -6186 424338
rect -6806 388658 -6774 388894
rect -6538 388658 -6454 388894
rect -6218 388658 -6186 388894
rect -6806 388574 -6186 388658
rect -6806 388338 -6774 388574
rect -6538 388338 -6454 388574
rect -6218 388338 -6186 388574
rect -6806 352894 -6186 388338
rect -6806 352658 -6774 352894
rect -6538 352658 -6454 352894
rect -6218 352658 -6186 352894
rect -6806 352574 -6186 352658
rect -6806 352338 -6774 352574
rect -6538 352338 -6454 352574
rect -6218 352338 -6186 352574
rect -6806 316894 -6186 352338
rect -6806 316658 -6774 316894
rect -6538 316658 -6454 316894
rect -6218 316658 -6186 316894
rect -6806 316574 -6186 316658
rect -6806 316338 -6774 316574
rect -6538 316338 -6454 316574
rect -6218 316338 -6186 316574
rect -6806 280894 -6186 316338
rect -6806 280658 -6774 280894
rect -6538 280658 -6454 280894
rect -6218 280658 -6186 280894
rect -6806 280574 -6186 280658
rect -6806 280338 -6774 280574
rect -6538 280338 -6454 280574
rect -6218 280338 -6186 280574
rect -6806 244894 -6186 280338
rect -6806 244658 -6774 244894
rect -6538 244658 -6454 244894
rect -6218 244658 -6186 244894
rect -6806 244574 -6186 244658
rect -6806 244338 -6774 244574
rect -6538 244338 -6454 244574
rect -6218 244338 -6186 244574
rect -6806 208894 -6186 244338
rect -6806 208658 -6774 208894
rect -6538 208658 -6454 208894
rect -6218 208658 -6186 208894
rect -6806 208574 -6186 208658
rect -6806 208338 -6774 208574
rect -6538 208338 -6454 208574
rect -6218 208338 -6186 208574
rect -6806 172894 -6186 208338
rect -6806 172658 -6774 172894
rect -6538 172658 -6454 172894
rect -6218 172658 -6186 172894
rect -6806 172574 -6186 172658
rect -6806 172338 -6774 172574
rect -6538 172338 -6454 172574
rect -6218 172338 -6186 172574
rect -6806 136894 -6186 172338
rect -6806 136658 -6774 136894
rect -6538 136658 -6454 136894
rect -6218 136658 -6186 136894
rect -6806 136574 -6186 136658
rect -6806 136338 -6774 136574
rect -6538 136338 -6454 136574
rect -6218 136338 -6186 136574
rect -6806 100894 -6186 136338
rect -6806 100658 -6774 100894
rect -6538 100658 -6454 100894
rect -6218 100658 -6186 100894
rect -6806 100574 -6186 100658
rect -6806 100338 -6774 100574
rect -6538 100338 -6454 100574
rect -6218 100338 -6186 100574
rect -6806 64894 -6186 100338
rect -6806 64658 -6774 64894
rect -6538 64658 -6454 64894
rect -6218 64658 -6186 64894
rect -6806 64574 -6186 64658
rect -6806 64338 -6774 64574
rect -6538 64338 -6454 64574
rect -6218 64338 -6186 64574
rect -6806 28894 -6186 64338
rect -6806 28658 -6774 28894
rect -6538 28658 -6454 28894
rect -6218 28658 -6186 28894
rect -6806 28574 -6186 28658
rect -6806 28338 -6774 28574
rect -6538 28338 -6454 28574
rect -6218 28338 -6186 28574
rect -6806 -5146 -6186 28338
rect -5846 708678 -5226 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 -5226 708678
rect -5846 708358 -5226 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 -5226 708358
rect -5846 694894 -5226 708122
rect 9234 708678 9854 709670
rect 9234 708442 9266 708678
rect 9502 708442 9586 708678
rect 9822 708442 9854 708678
rect 9234 708358 9854 708442
rect 9234 708122 9266 708358
rect 9502 708122 9586 708358
rect 9822 708122 9854 708358
rect -5846 694658 -5814 694894
rect -5578 694658 -5494 694894
rect -5258 694658 -5226 694894
rect -5846 694574 -5226 694658
rect -5846 694338 -5814 694574
rect -5578 694338 -5494 694574
rect -5258 694338 -5226 694574
rect -5846 658894 -5226 694338
rect -5846 658658 -5814 658894
rect -5578 658658 -5494 658894
rect -5258 658658 -5226 658894
rect -5846 658574 -5226 658658
rect -5846 658338 -5814 658574
rect -5578 658338 -5494 658574
rect -5258 658338 -5226 658574
rect -5846 622894 -5226 658338
rect -5846 622658 -5814 622894
rect -5578 622658 -5494 622894
rect -5258 622658 -5226 622894
rect -5846 622574 -5226 622658
rect -5846 622338 -5814 622574
rect -5578 622338 -5494 622574
rect -5258 622338 -5226 622574
rect -5846 586894 -5226 622338
rect -5846 586658 -5814 586894
rect -5578 586658 -5494 586894
rect -5258 586658 -5226 586894
rect -5846 586574 -5226 586658
rect -5846 586338 -5814 586574
rect -5578 586338 -5494 586574
rect -5258 586338 -5226 586574
rect -5846 550894 -5226 586338
rect -5846 550658 -5814 550894
rect -5578 550658 -5494 550894
rect -5258 550658 -5226 550894
rect -5846 550574 -5226 550658
rect -5846 550338 -5814 550574
rect -5578 550338 -5494 550574
rect -5258 550338 -5226 550574
rect -5846 514894 -5226 550338
rect -5846 514658 -5814 514894
rect -5578 514658 -5494 514894
rect -5258 514658 -5226 514894
rect -5846 514574 -5226 514658
rect -5846 514338 -5814 514574
rect -5578 514338 -5494 514574
rect -5258 514338 -5226 514574
rect -5846 478894 -5226 514338
rect -5846 478658 -5814 478894
rect -5578 478658 -5494 478894
rect -5258 478658 -5226 478894
rect -5846 478574 -5226 478658
rect -5846 478338 -5814 478574
rect -5578 478338 -5494 478574
rect -5258 478338 -5226 478574
rect -5846 442894 -5226 478338
rect -5846 442658 -5814 442894
rect -5578 442658 -5494 442894
rect -5258 442658 -5226 442894
rect -5846 442574 -5226 442658
rect -5846 442338 -5814 442574
rect -5578 442338 -5494 442574
rect -5258 442338 -5226 442574
rect -5846 406894 -5226 442338
rect -5846 406658 -5814 406894
rect -5578 406658 -5494 406894
rect -5258 406658 -5226 406894
rect -5846 406574 -5226 406658
rect -5846 406338 -5814 406574
rect -5578 406338 -5494 406574
rect -5258 406338 -5226 406574
rect -5846 370894 -5226 406338
rect -5846 370658 -5814 370894
rect -5578 370658 -5494 370894
rect -5258 370658 -5226 370894
rect -5846 370574 -5226 370658
rect -5846 370338 -5814 370574
rect -5578 370338 -5494 370574
rect -5258 370338 -5226 370574
rect -5846 334894 -5226 370338
rect -5846 334658 -5814 334894
rect -5578 334658 -5494 334894
rect -5258 334658 -5226 334894
rect -5846 334574 -5226 334658
rect -5846 334338 -5814 334574
rect -5578 334338 -5494 334574
rect -5258 334338 -5226 334574
rect -5846 298894 -5226 334338
rect -5846 298658 -5814 298894
rect -5578 298658 -5494 298894
rect -5258 298658 -5226 298894
rect -5846 298574 -5226 298658
rect -5846 298338 -5814 298574
rect -5578 298338 -5494 298574
rect -5258 298338 -5226 298574
rect -5846 262894 -5226 298338
rect -5846 262658 -5814 262894
rect -5578 262658 -5494 262894
rect -5258 262658 -5226 262894
rect -5846 262574 -5226 262658
rect -5846 262338 -5814 262574
rect -5578 262338 -5494 262574
rect -5258 262338 -5226 262574
rect -5846 226894 -5226 262338
rect -5846 226658 -5814 226894
rect -5578 226658 -5494 226894
rect -5258 226658 -5226 226894
rect -5846 226574 -5226 226658
rect -5846 226338 -5814 226574
rect -5578 226338 -5494 226574
rect -5258 226338 -5226 226574
rect -5846 190894 -5226 226338
rect -5846 190658 -5814 190894
rect -5578 190658 -5494 190894
rect -5258 190658 -5226 190894
rect -5846 190574 -5226 190658
rect -5846 190338 -5814 190574
rect -5578 190338 -5494 190574
rect -5258 190338 -5226 190574
rect -5846 154894 -5226 190338
rect -5846 154658 -5814 154894
rect -5578 154658 -5494 154894
rect -5258 154658 -5226 154894
rect -5846 154574 -5226 154658
rect -5846 154338 -5814 154574
rect -5578 154338 -5494 154574
rect -5258 154338 -5226 154574
rect -5846 118894 -5226 154338
rect -5846 118658 -5814 118894
rect -5578 118658 -5494 118894
rect -5258 118658 -5226 118894
rect -5846 118574 -5226 118658
rect -5846 118338 -5814 118574
rect -5578 118338 -5494 118574
rect -5258 118338 -5226 118574
rect -5846 82894 -5226 118338
rect -5846 82658 -5814 82894
rect -5578 82658 -5494 82894
rect -5258 82658 -5226 82894
rect -5846 82574 -5226 82658
rect -5846 82338 -5814 82574
rect -5578 82338 -5494 82574
rect -5258 82338 -5226 82574
rect -5846 46894 -5226 82338
rect -5846 46658 -5814 46894
rect -5578 46658 -5494 46894
rect -5258 46658 -5226 46894
rect -5846 46574 -5226 46658
rect -5846 46338 -5814 46574
rect -5578 46338 -5494 46574
rect -5258 46338 -5226 46574
rect -5846 10894 -5226 46338
rect -5846 10658 -5814 10894
rect -5578 10658 -5494 10894
rect -5258 10658 -5226 10894
rect -5846 10574 -5226 10658
rect -5846 10338 -5814 10574
rect -5578 10338 -5494 10574
rect -5258 10338 -5226 10574
rect -5846 -4186 -5226 10338
rect -4886 707718 -4266 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 -4266 707718
rect -4886 707398 -4266 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 -4266 707398
rect -4886 673174 -4266 707162
rect -4886 672938 -4854 673174
rect -4618 672938 -4534 673174
rect -4298 672938 -4266 673174
rect -4886 672854 -4266 672938
rect -4886 672618 -4854 672854
rect -4618 672618 -4534 672854
rect -4298 672618 -4266 672854
rect -4886 637174 -4266 672618
rect -4886 636938 -4854 637174
rect -4618 636938 -4534 637174
rect -4298 636938 -4266 637174
rect -4886 636854 -4266 636938
rect -4886 636618 -4854 636854
rect -4618 636618 -4534 636854
rect -4298 636618 -4266 636854
rect -4886 601174 -4266 636618
rect -4886 600938 -4854 601174
rect -4618 600938 -4534 601174
rect -4298 600938 -4266 601174
rect -4886 600854 -4266 600938
rect -4886 600618 -4854 600854
rect -4618 600618 -4534 600854
rect -4298 600618 -4266 600854
rect -4886 565174 -4266 600618
rect -4886 564938 -4854 565174
rect -4618 564938 -4534 565174
rect -4298 564938 -4266 565174
rect -4886 564854 -4266 564938
rect -4886 564618 -4854 564854
rect -4618 564618 -4534 564854
rect -4298 564618 -4266 564854
rect -4886 529174 -4266 564618
rect -4886 528938 -4854 529174
rect -4618 528938 -4534 529174
rect -4298 528938 -4266 529174
rect -4886 528854 -4266 528938
rect -4886 528618 -4854 528854
rect -4618 528618 -4534 528854
rect -4298 528618 -4266 528854
rect -4886 493174 -4266 528618
rect -4886 492938 -4854 493174
rect -4618 492938 -4534 493174
rect -4298 492938 -4266 493174
rect -4886 492854 -4266 492938
rect -4886 492618 -4854 492854
rect -4618 492618 -4534 492854
rect -4298 492618 -4266 492854
rect -4886 457174 -4266 492618
rect -4886 456938 -4854 457174
rect -4618 456938 -4534 457174
rect -4298 456938 -4266 457174
rect -4886 456854 -4266 456938
rect -4886 456618 -4854 456854
rect -4618 456618 -4534 456854
rect -4298 456618 -4266 456854
rect -4886 421174 -4266 456618
rect -4886 420938 -4854 421174
rect -4618 420938 -4534 421174
rect -4298 420938 -4266 421174
rect -4886 420854 -4266 420938
rect -4886 420618 -4854 420854
rect -4618 420618 -4534 420854
rect -4298 420618 -4266 420854
rect -4886 385174 -4266 420618
rect -4886 384938 -4854 385174
rect -4618 384938 -4534 385174
rect -4298 384938 -4266 385174
rect -4886 384854 -4266 384938
rect -4886 384618 -4854 384854
rect -4618 384618 -4534 384854
rect -4298 384618 -4266 384854
rect -4886 349174 -4266 384618
rect -4886 348938 -4854 349174
rect -4618 348938 -4534 349174
rect -4298 348938 -4266 349174
rect -4886 348854 -4266 348938
rect -4886 348618 -4854 348854
rect -4618 348618 -4534 348854
rect -4298 348618 -4266 348854
rect -4886 313174 -4266 348618
rect -4886 312938 -4854 313174
rect -4618 312938 -4534 313174
rect -4298 312938 -4266 313174
rect -4886 312854 -4266 312938
rect -4886 312618 -4854 312854
rect -4618 312618 -4534 312854
rect -4298 312618 -4266 312854
rect -4886 277174 -4266 312618
rect -4886 276938 -4854 277174
rect -4618 276938 -4534 277174
rect -4298 276938 -4266 277174
rect -4886 276854 -4266 276938
rect -4886 276618 -4854 276854
rect -4618 276618 -4534 276854
rect -4298 276618 -4266 276854
rect -4886 241174 -4266 276618
rect -4886 240938 -4854 241174
rect -4618 240938 -4534 241174
rect -4298 240938 -4266 241174
rect -4886 240854 -4266 240938
rect -4886 240618 -4854 240854
rect -4618 240618 -4534 240854
rect -4298 240618 -4266 240854
rect -4886 205174 -4266 240618
rect -4886 204938 -4854 205174
rect -4618 204938 -4534 205174
rect -4298 204938 -4266 205174
rect -4886 204854 -4266 204938
rect -4886 204618 -4854 204854
rect -4618 204618 -4534 204854
rect -4298 204618 -4266 204854
rect -4886 169174 -4266 204618
rect -4886 168938 -4854 169174
rect -4618 168938 -4534 169174
rect -4298 168938 -4266 169174
rect -4886 168854 -4266 168938
rect -4886 168618 -4854 168854
rect -4618 168618 -4534 168854
rect -4298 168618 -4266 168854
rect -4886 133174 -4266 168618
rect -4886 132938 -4854 133174
rect -4618 132938 -4534 133174
rect -4298 132938 -4266 133174
rect -4886 132854 -4266 132938
rect -4886 132618 -4854 132854
rect -4618 132618 -4534 132854
rect -4298 132618 -4266 132854
rect -4886 97174 -4266 132618
rect -4886 96938 -4854 97174
rect -4618 96938 -4534 97174
rect -4298 96938 -4266 97174
rect -4886 96854 -4266 96938
rect -4886 96618 -4854 96854
rect -4618 96618 -4534 96854
rect -4298 96618 -4266 96854
rect -4886 61174 -4266 96618
rect -4886 60938 -4854 61174
rect -4618 60938 -4534 61174
rect -4298 60938 -4266 61174
rect -4886 60854 -4266 60938
rect -4886 60618 -4854 60854
rect -4618 60618 -4534 60854
rect -4298 60618 -4266 60854
rect -4886 25174 -4266 60618
rect -4886 24938 -4854 25174
rect -4618 24938 -4534 25174
rect -4298 24938 -4266 25174
rect -4886 24854 -4266 24938
rect -4886 24618 -4854 24854
rect -4618 24618 -4534 24854
rect -4298 24618 -4266 24854
rect -4886 -3226 -4266 24618
rect -3926 706758 -3306 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 -3306 706758
rect -3926 706438 -3306 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 -3306 706438
rect -3926 691174 -3306 706202
rect 5514 706758 6134 707750
rect 5514 706522 5546 706758
rect 5782 706522 5866 706758
rect 6102 706522 6134 706758
rect 5514 706438 6134 706522
rect 5514 706202 5546 706438
rect 5782 706202 5866 706438
rect 6102 706202 6134 706438
rect -3926 690938 -3894 691174
rect -3658 690938 -3574 691174
rect -3338 690938 -3306 691174
rect -3926 690854 -3306 690938
rect -3926 690618 -3894 690854
rect -3658 690618 -3574 690854
rect -3338 690618 -3306 690854
rect -3926 655174 -3306 690618
rect -3926 654938 -3894 655174
rect -3658 654938 -3574 655174
rect -3338 654938 -3306 655174
rect -3926 654854 -3306 654938
rect -3926 654618 -3894 654854
rect -3658 654618 -3574 654854
rect -3338 654618 -3306 654854
rect -3926 619174 -3306 654618
rect -3926 618938 -3894 619174
rect -3658 618938 -3574 619174
rect -3338 618938 -3306 619174
rect -3926 618854 -3306 618938
rect -3926 618618 -3894 618854
rect -3658 618618 -3574 618854
rect -3338 618618 -3306 618854
rect -3926 583174 -3306 618618
rect -3926 582938 -3894 583174
rect -3658 582938 -3574 583174
rect -3338 582938 -3306 583174
rect -3926 582854 -3306 582938
rect -3926 582618 -3894 582854
rect -3658 582618 -3574 582854
rect -3338 582618 -3306 582854
rect -3926 547174 -3306 582618
rect -3926 546938 -3894 547174
rect -3658 546938 -3574 547174
rect -3338 546938 -3306 547174
rect -3926 546854 -3306 546938
rect -3926 546618 -3894 546854
rect -3658 546618 -3574 546854
rect -3338 546618 -3306 546854
rect -3926 511174 -3306 546618
rect -3926 510938 -3894 511174
rect -3658 510938 -3574 511174
rect -3338 510938 -3306 511174
rect -3926 510854 -3306 510938
rect -3926 510618 -3894 510854
rect -3658 510618 -3574 510854
rect -3338 510618 -3306 510854
rect -3926 475174 -3306 510618
rect -3926 474938 -3894 475174
rect -3658 474938 -3574 475174
rect -3338 474938 -3306 475174
rect -3926 474854 -3306 474938
rect -3926 474618 -3894 474854
rect -3658 474618 -3574 474854
rect -3338 474618 -3306 474854
rect -3926 439174 -3306 474618
rect -3926 438938 -3894 439174
rect -3658 438938 -3574 439174
rect -3338 438938 -3306 439174
rect -3926 438854 -3306 438938
rect -3926 438618 -3894 438854
rect -3658 438618 -3574 438854
rect -3338 438618 -3306 438854
rect -3926 403174 -3306 438618
rect -3926 402938 -3894 403174
rect -3658 402938 -3574 403174
rect -3338 402938 -3306 403174
rect -3926 402854 -3306 402938
rect -3926 402618 -3894 402854
rect -3658 402618 -3574 402854
rect -3338 402618 -3306 402854
rect -3926 367174 -3306 402618
rect -3926 366938 -3894 367174
rect -3658 366938 -3574 367174
rect -3338 366938 -3306 367174
rect -3926 366854 -3306 366938
rect -3926 366618 -3894 366854
rect -3658 366618 -3574 366854
rect -3338 366618 -3306 366854
rect -3926 331174 -3306 366618
rect -3926 330938 -3894 331174
rect -3658 330938 -3574 331174
rect -3338 330938 -3306 331174
rect -3926 330854 -3306 330938
rect -3926 330618 -3894 330854
rect -3658 330618 -3574 330854
rect -3338 330618 -3306 330854
rect -3926 295174 -3306 330618
rect -3926 294938 -3894 295174
rect -3658 294938 -3574 295174
rect -3338 294938 -3306 295174
rect -3926 294854 -3306 294938
rect -3926 294618 -3894 294854
rect -3658 294618 -3574 294854
rect -3338 294618 -3306 294854
rect -3926 259174 -3306 294618
rect -3926 258938 -3894 259174
rect -3658 258938 -3574 259174
rect -3338 258938 -3306 259174
rect -3926 258854 -3306 258938
rect -3926 258618 -3894 258854
rect -3658 258618 -3574 258854
rect -3338 258618 -3306 258854
rect -3926 223174 -3306 258618
rect -3926 222938 -3894 223174
rect -3658 222938 -3574 223174
rect -3338 222938 -3306 223174
rect -3926 222854 -3306 222938
rect -3926 222618 -3894 222854
rect -3658 222618 -3574 222854
rect -3338 222618 -3306 222854
rect -3926 187174 -3306 222618
rect -3926 186938 -3894 187174
rect -3658 186938 -3574 187174
rect -3338 186938 -3306 187174
rect -3926 186854 -3306 186938
rect -3926 186618 -3894 186854
rect -3658 186618 -3574 186854
rect -3338 186618 -3306 186854
rect -3926 151174 -3306 186618
rect -3926 150938 -3894 151174
rect -3658 150938 -3574 151174
rect -3338 150938 -3306 151174
rect -3926 150854 -3306 150938
rect -3926 150618 -3894 150854
rect -3658 150618 -3574 150854
rect -3338 150618 -3306 150854
rect -3926 115174 -3306 150618
rect -3926 114938 -3894 115174
rect -3658 114938 -3574 115174
rect -3338 114938 -3306 115174
rect -3926 114854 -3306 114938
rect -3926 114618 -3894 114854
rect -3658 114618 -3574 114854
rect -3338 114618 -3306 114854
rect -3926 79174 -3306 114618
rect -3926 78938 -3894 79174
rect -3658 78938 -3574 79174
rect -3338 78938 -3306 79174
rect -3926 78854 -3306 78938
rect -3926 78618 -3894 78854
rect -3658 78618 -3574 78854
rect -3338 78618 -3306 78854
rect -3926 43174 -3306 78618
rect -3926 42938 -3894 43174
rect -3658 42938 -3574 43174
rect -3338 42938 -3306 43174
rect -3926 42854 -3306 42938
rect -3926 42618 -3894 42854
rect -3658 42618 -3574 42854
rect -3338 42618 -3306 42854
rect -3926 7174 -3306 42618
rect -3926 6938 -3894 7174
rect -3658 6938 -3574 7174
rect -3338 6938 -3306 7174
rect -3926 6854 -3306 6938
rect -3926 6618 -3894 6854
rect -3658 6618 -3574 6854
rect -3338 6618 -3306 6854
rect -3926 -2266 -3306 6618
rect -2966 705798 -2346 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 -2346 705798
rect -2966 705478 -2346 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 -2346 705478
rect -2966 669454 -2346 705242
rect -2966 669218 -2934 669454
rect -2698 669218 -2614 669454
rect -2378 669218 -2346 669454
rect -2966 669134 -2346 669218
rect -2966 668898 -2934 669134
rect -2698 668898 -2614 669134
rect -2378 668898 -2346 669134
rect -2966 633454 -2346 668898
rect -2966 633218 -2934 633454
rect -2698 633218 -2614 633454
rect -2378 633218 -2346 633454
rect -2966 633134 -2346 633218
rect -2966 632898 -2934 633134
rect -2698 632898 -2614 633134
rect -2378 632898 -2346 633134
rect -2966 597454 -2346 632898
rect -2966 597218 -2934 597454
rect -2698 597218 -2614 597454
rect -2378 597218 -2346 597454
rect -2966 597134 -2346 597218
rect -2966 596898 -2934 597134
rect -2698 596898 -2614 597134
rect -2378 596898 -2346 597134
rect -2966 561454 -2346 596898
rect -2966 561218 -2934 561454
rect -2698 561218 -2614 561454
rect -2378 561218 -2346 561454
rect -2966 561134 -2346 561218
rect -2966 560898 -2934 561134
rect -2698 560898 -2614 561134
rect -2378 560898 -2346 561134
rect -2966 525454 -2346 560898
rect -2966 525218 -2934 525454
rect -2698 525218 -2614 525454
rect -2378 525218 -2346 525454
rect -2966 525134 -2346 525218
rect -2966 524898 -2934 525134
rect -2698 524898 -2614 525134
rect -2378 524898 -2346 525134
rect -2966 489454 -2346 524898
rect -2966 489218 -2934 489454
rect -2698 489218 -2614 489454
rect -2378 489218 -2346 489454
rect -2966 489134 -2346 489218
rect -2966 488898 -2934 489134
rect -2698 488898 -2614 489134
rect -2378 488898 -2346 489134
rect -2966 453454 -2346 488898
rect -2966 453218 -2934 453454
rect -2698 453218 -2614 453454
rect -2378 453218 -2346 453454
rect -2966 453134 -2346 453218
rect -2966 452898 -2934 453134
rect -2698 452898 -2614 453134
rect -2378 452898 -2346 453134
rect -2966 417454 -2346 452898
rect -2966 417218 -2934 417454
rect -2698 417218 -2614 417454
rect -2378 417218 -2346 417454
rect -2966 417134 -2346 417218
rect -2966 416898 -2934 417134
rect -2698 416898 -2614 417134
rect -2378 416898 -2346 417134
rect -2966 381454 -2346 416898
rect -2966 381218 -2934 381454
rect -2698 381218 -2614 381454
rect -2378 381218 -2346 381454
rect -2966 381134 -2346 381218
rect -2966 380898 -2934 381134
rect -2698 380898 -2614 381134
rect -2378 380898 -2346 381134
rect -2966 345454 -2346 380898
rect -2966 345218 -2934 345454
rect -2698 345218 -2614 345454
rect -2378 345218 -2346 345454
rect -2966 345134 -2346 345218
rect -2966 344898 -2934 345134
rect -2698 344898 -2614 345134
rect -2378 344898 -2346 345134
rect -2966 309454 -2346 344898
rect -2966 309218 -2934 309454
rect -2698 309218 -2614 309454
rect -2378 309218 -2346 309454
rect -2966 309134 -2346 309218
rect -2966 308898 -2934 309134
rect -2698 308898 -2614 309134
rect -2378 308898 -2346 309134
rect -2966 273454 -2346 308898
rect -2966 273218 -2934 273454
rect -2698 273218 -2614 273454
rect -2378 273218 -2346 273454
rect -2966 273134 -2346 273218
rect -2966 272898 -2934 273134
rect -2698 272898 -2614 273134
rect -2378 272898 -2346 273134
rect -2966 237454 -2346 272898
rect -2966 237218 -2934 237454
rect -2698 237218 -2614 237454
rect -2378 237218 -2346 237454
rect -2966 237134 -2346 237218
rect -2966 236898 -2934 237134
rect -2698 236898 -2614 237134
rect -2378 236898 -2346 237134
rect -2966 201454 -2346 236898
rect -2966 201218 -2934 201454
rect -2698 201218 -2614 201454
rect -2378 201218 -2346 201454
rect -2966 201134 -2346 201218
rect -2966 200898 -2934 201134
rect -2698 200898 -2614 201134
rect -2378 200898 -2346 201134
rect -2966 165454 -2346 200898
rect -2966 165218 -2934 165454
rect -2698 165218 -2614 165454
rect -2378 165218 -2346 165454
rect -2966 165134 -2346 165218
rect -2966 164898 -2934 165134
rect -2698 164898 -2614 165134
rect -2378 164898 -2346 165134
rect -2966 129454 -2346 164898
rect -2966 129218 -2934 129454
rect -2698 129218 -2614 129454
rect -2378 129218 -2346 129454
rect -2966 129134 -2346 129218
rect -2966 128898 -2934 129134
rect -2698 128898 -2614 129134
rect -2378 128898 -2346 129134
rect -2966 93454 -2346 128898
rect -2966 93218 -2934 93454
rect -2698 93218 -2614 93454
rect -2378 93218 -2346 93454
rect -2966 93134 -2346 93218
rect -2966 92898 -2934 93134
rect -2698 92898 -2614 93134
rect -2378 92898 -2346 93134
rect -2966 57454 -2346 92898
rect -2966 57218 -2934 57454
rect -2698 57218 -2614 57454
rect -2378 57218 -2346 57454
rect -2966 57134 -2346 57218
rect -2966 56898 -2934 57134
rect -2698 56898 -2614 57134
rect -2378 56898 -2346 57134
rect -2966 21454 -2346 56898
rect -2966 21218 -2934 21454
rect -2698 21218 -2614 21454
rect -2378 21218 -2346 21454
rect -2966 21134 -2346 21218
rect -2966 20898 -2934 21134
rect -2698 20898 -2614 21134
rect -2378 20898 -2346 21134
rect -2966 -1306 -2346 20898
rect -2006 704838 -1386 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 -1386 704838
rect -2006 704518 -1386 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 -1386 704518
rect -2006 687454 -1386 704282
rect -2006 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 -1386 687454
rect -2006 687134 -1386 687218
rect -2006 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 -1386 687134
rect -2006 651454 -1386 686898
rect -2006 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 -1386 651454
rect -2006 651134 -1386 651218
rect -2006 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 -1386 651134
rect -2006 615454 -1386 650898
rect -2006 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 -1386 615454
rect -2006 615134 -1386 615218
rect -2006 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 -1386 615134
rect -2006 579454 -1386 614898
rect -2006 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 -1386 579454
rect -2006 579134 -1386 579218
rect -2006 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 -1386 579134
rect -2006 543454 -1386 578898
rect -2006 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 -1386 543454
rect -2006 543134 -1386 543218
rect -2006 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 -1386 543134
rect -2006 507454 -1386 542898
rect -2006 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 -1386 507454
rect -2006 507134 -1386 507218
rect -2006 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 -1386 507134
rect -2006 471454 -1386 506898
rect -2006 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 -1386 471454
rect -2006 471134 -1386 471218
rect -2006 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 -1386 471134
rect -2006 435454 -1386 470898
rect -2006 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 -1386 435454
rect -2006 435134 -1386 435218
rect -2006 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 -1386 435134
rect -2006 399454 -1386 434898
rect -2006 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 -1386 399454
rect -2006 399134 -1386 399218
rect -2006 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 -1386 399134
rect -2006 363454 -1386 398898
rect -2006 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 -1386 363454
rect -2006 363134 -1386 363218
rect -2006 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 -1386 363134
rect -2006 327454 -1386 362898
rect -2006 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 -1386 327454
rect -2006 327134 -1386 327218
rect -2006 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 -1386 327134
rect -2006 291454 -1386 326898
rect -2006 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 -1386 291454
rect -2006 291134 -1386 291218
rect -2006 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 -1386 291134
rect -2006 255454 -1386 290898
rect -2006 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 -1386 255454
rect -2006 255134 -1386 255218
rect -2006 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 -1386 255134
rect -2006 219454 -1386 254898
rect -2006 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 -1386 219454
rect -2006 219134 -1386 219218
rect -2006 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 -1386 219134
rect -2006 183454 -1386 218898
rect -2006 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 -1386 183454
rect -2006 183134 -1386 183218
rect -2006 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 -1386 183134
rect -2006 147454 -1386 182898
rect -2006 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 -1386 147454
rect -2006 147134 -1386 147218
rect -2006 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 -1386 147134
rect -2006 111454 -1386 146898
rect -2006 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 -1386 111454
rect -2006 111134 -1386 111218
rect -2006 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 -1386 111134
rect -2006 75454 -1386 110898
rect -2006 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 -1386 75454
rect -2006 75134 -1386 75218
rect -2006 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 -1386 75134
rect -2006 39454 -1386 74898
rect -2006 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 -1386 39454
rect -2006 39134 -1386 39218
rect -2006 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 -1386 39134
rect -2006 3454 -1386 38898
rect -2006 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 -1386 3454
rect -2006 3134 -1386 3218
rect -2006 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 -1386 3134
rect -2006 -346 -1386 2898
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 -1386 -346
rect -2006 -666 -1386 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 -1386 -666
rect -2006 -934 -1386 -902
rect 1794 704838 2414 705830
rect 1794 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 2414 704838
rect 1794 704518 2414 704602
rect 1794 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 2414 704518
rect 1794 687454 2414 704282
rect 1794 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 2414 687454
rect 1794 687134 2414 687218
rect 1794 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 2414 687134
rect 1794 651454 2414 686898
rect 1794 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 2414 651454
rect 1794 651134 2414 651218
rect 1794 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 2414 651134
rect 1794 615454 2414 650898
rect 1794 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 2414 615454
rect 1794 615134 2414 615218
rect 1794 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 2414 615134
rect 1794 579454 2414 614898
rect 1794 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 2414 579454
rect 1794 579134 2414 579218
rect 1794 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 2414 579134
rect 1794 543454 2414 578898
rect 1794 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 2414 543454
rect 1794 543134 2414 543218
rect 1794 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 2414 543134
rect 1794 507454 2414 542898
rect 1794 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 2414 507454
rect 1794 507134 2414 507218
rect 1794 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 2414 507134
rect 1794 471454 2414 506898
rect 1794 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 2414 471454
rect 1794 471134 2414 471218
rect 1794 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 2414 471134
rect 1794 435454 2414 470898
rect 1794 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 2414 435454
rect 1794 435134 2414 435218
rect 1794 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 2414 435134
rect 1794 399454 2414 434898
rect 1794 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 2414 399454
rect 1794 399134 2414 399218
rect 1794 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 2414 399134
rect 1794 363454 2414 398898
rect 1794 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 2414 363454
rect 1794 363134 2414 363218
rect 1794 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 2414 363134
rect 1794 327454 2414 362898
rect 1794 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 2414 327454
rect 1794 327134 2414 327218
rect 1794 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 2414 327134
rect 1794 291454 2414 326898
rect 1794 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 2414 291454
rect 1794 291134 2414 291218
rect 1794 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 2414 291134
rect 1794 255454 2414 290898
rect 1794 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 2414 255454
rect 1794 255134 2414 255218
rect 1794 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 2414 255134
rect 1794 219454 2414 254898
rect 1794 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 2414 219454
rect 1794 219134 2414 219218
rect 1794 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 2414 219134
rect 1794 183454 2414 218898
rect 1794 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 2414 183454
rect 1794 183134 2414 183218
rect 1794 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 2414 183134
rect 1794 147454 2414 182898
rect 1794 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 2414 147454
rect 1794 147134 2414 147218
rect 1794 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 2414 147134
rect 1794 111454 2414 146898
rect 1794 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 2414 111454
rect 1794 111134 2414 111218
rect 1794 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 2414 111134
rect 1794 75454 2414 110898
rect 1794 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 2414 75454
rect 1794 75134 2414 75218
rect 1794 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 2414 75134
rect 1794 39454 2414 74898
rect 1794 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 2414 39454
rect 1794 39134 2414 39218
rect 1794 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 2414 39134
rect 1794 3454 2414 38898
rect 1794 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 2414 3454
rect 1794 3134 2414 3218
rect 1794 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 2414 3134
rect 1794 -346 2414 2898
rect 1794 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 2414 -346
rect 1794 -666 2414 -582
rect 1794 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 2414 -666
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 -2346 -1306
rect -2966 -1626 -2346 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 -2346 -1626
rect -2966 -1894 -2346 -1862
rect 1794 -1894 2414 -902
rect 5514 691174 6134 706202
rect 5514 690938 5546 691174
rect 5782 690938 5866 691174
rect 6102 690938 6134 691174
rect 5514 690854 6134 690938
rect 5514 690618 5546 690854
rect 5782 690618 5866 690854
rect 6102 690618 6134 690854
rect 5514 655174 6134 690618
rect 5514 654938 5546 655174
rect 5782 654938 5866 655174
rect 6102 654938 6134 655174
rect 5514 654854 6134 654938
rect 5514 654618 5546 654854
rect 5782 654618 5866 654854
rect 6102 654618 6134 654854
rect 5514 619174 6134 654618
rect 5514 618938 5546 619174
rect 5782 618938 5866 619174
rect 6102 618938 6134 619174
rect 5514 618854 6134 618938
rect 5514 618618 5546 618854
rect 5782 618618 5866 618854
rect 6102 618618 6134 618854
rect 5514 583174 6134 618618
rect 5514 582938 5546 583174
rect 5782 582938 5866 583174
rect 6102 582938 6134 583174
rect 5514 582854 6134 582938
rect 5514 582618 5546 582854
rect 5782 582618 5866 582854
rect 6102 582618 6134 582854
rect 5514 547174 6134 582618
rect 5514 546938 5546 547174
rect 5782 546938 5866 547174
rect 6102 546938 6134 547174
rect 5514 546854 6134 546938
rect 5514 546618 5546 546854
rect 5782 546618 5866 546854
rect 6102 546618 6134 546854
rect 5514 511174 6134 546618
rect 5514 510938 5546 511174
rect 5782 510938 5866 511174
rect 6102 510938 6134 511174
rect 5514 510854 6134 510938
rect 5514 510618 5546 510854
rect 5782 510618 5866 510854
rect 6102 510618 6134 510854
rect 5514 475174 6134 510618
rect 5514 474938 5546 475174
rect 5782 474938 5866 475174
rect 6102 474938 6134 475174
rect 5514 474854 6134 474938
rect 5514 474618 5546 474854
rect 5782 474618 5866 474854
rect 6102 474618 6134 474854
rect 5514 439174 6134 474618
rect 5514 438938 5546 439174
rect 5782 438938 5866 439174
rect 6102 438938 6134 439174
rect 5514 438854 6134 438938
rect 5514 438618 5546 438854
rect 5782 438618 5866 438854
rect 6102 438618 6134 438854
rect 5514 403174 6134 438618
rect 5514 402938 5546 403174
rect 5782 402938 5866 403174
rect 6102 402938 6134 403174
rect 5514 402854 6134 402938
rect 5514 402618 5546 402854
rect 5782 402618 5866 402854
rect 6102 402618 6134 402854
rect 5514 367174 6134 402618
rect 5514 366938 5546 367174
rect 5782 366938 5866 367174
rect 6102 366938 6134 367174
rect 5514 366854 6134 366938
rect 5514 366618 5546 366854
rect 5782 366618 5866 366854
rect 6102 366618 6134 366854
rect 5514 331174 6134 366618
rect 5514 330938 5546 331174
rect 5782 330938 5866 331174
rect 6102 330938 6134 331174
rect 5514 330854 6134 330938
rect 5514 330618 5546 330854
rect 5782 330618 5866 330854
rect 6102 330618 6134 330854
rect 5514 295174 6134 330618
rect 5514 294938 5546 295174
rect 5782 294938 5866 295174
rect 6102 294938 6134 295174
rect 5514 294854 6134 294938
rect 5514 294618 5546 294854
rect 5782 294618 5866 294854
rect 6102 294618 6134 294854
rect 5514 259174 6134 294618
rect 5514 258938 5546 259174
rect 5782 258938 5866 259174
rect 6102 258938 6134 259174
rect 5514 258854 6134 258938
rect 5514 258618 5546 258854
rect 5782 258618 5866 258854
rect 6102 258618 6134 258854
rect 5514 223174 6134 258618
rect 5514 222938 5546 223174
rect 5782 222938 5866 223174
rect 6102 222938 6134 223174
rect 5514 222854 6134 222938
rect 5514 222618 5546 222854
rect 5782 222618 5866 222854
rect 6102 222618 6134 222854
rect 5514 187174 6134 222618
rect 5514 186938 5546 187174
rect 5782 186938 5866 187174
rect 6102 186938 6134 187174
rect 5514 186854 6134 186938
rect 5514 186618 5546 186854
rect 5782 186618 5866 186854
rect 6102 186618 6134 186854
rect 5514 151174 6134 186618
rect 5514 150938 5546 151174
rect 5782 150938 5866 151174
rect 6102 150938 6134 151174
rect 5514 150854 6134 150938
rect 5514 150618 5546 150854
rect 5782 150618 5866 150854
rect 6102 150618 6134 150854
rect 5514 115174 6134 150618
rect 5514 114938 5546 115174
rect 5782 114938 5866 115174
rect 6102 114938 6134 115174
rect 5514 114854 6134 114938
rect 5514 114618 5546 114854
rect 5782 114618 5866 114854
rect 6102 114618 6134 114854
rect 5514 79174 6134 114618
rect 5514 78938 5546 79174
rect 5782 78938 5866 79174
rect 6102 78938 6134 79174
rect 5514 78854 6134 78938
rect 5514 78618 5546 78854
rect 5782 78618 5866 78854
rect 6102 78618 6134 78854
rect 5514 43174 6134 78618
rect 5514 42938 5546 43174
rect 5782 42938 5866 43174
rect 6102 42938 6134 43174
rect 5514 42854 6134 42938
rect 5514 42618 5546 42854
rect 5782 42618 5866 42854
rect 6102 42618 6134 42854
rect 5514 7174 6134 42618
rect 5514 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 6134 7174
rect 5514 6854 6134 6938
rect 5514 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 6134 6854
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 -3306 -2266
rect -3926 -2586 -3306 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 -3306 -2586
rect -3926 -2854 -3306 -2822
rect 5514 -2266 6134 6618
rect 5514 -2502 5546 -2266
rect 5782 -2502 5866 -2266
rect 6102 -2502 6134 -2266
rect 5514 -2586 6134 -2502
rect 5514 -2822 5546 -2586
rect 5782 -2822 5866 -2586
rect 6102 -2822 6134 -2586
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 -4266 -3226
rect -4886 -3546 -4266 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 -4266 -3546
rect -4886 -3814 -4266 -3782
rect 5514 -3814 6134 -2822
rect 9234 694894 9854 708122
rect 9234 694658 9266 694894
rect 9502 694658 9586 694894
rect 9822 694658 9854 694894
rect 9234 694574 9854 694658
rect 9234 694338 9266 694574
rect 9502 694338 9586 694574
rect 9822 694338 9854 694574
rect 9234 658894 9854 694338
rect 9234 658658 9266 658894
rect 9502 658658 9586 658894
rect 9822 658658 9854 658894
rect 9234 658574 9854 658658
rect 9234 658338 9266 658574
rect 9502 658338 9586 658574
rect 9822 658338 9854 658574
rect 9234 622894 9854 658338
rect 9234 622658 9266 622894
rect 9502 622658 9586 622894
rect 9822 622658 9854 622894
rect 9234 622574 9854 622658
rect 9234 622338 9266 622574
rect 9502 622338 9586 622574
rect 9822 622338 9854 622574
rect 9234 586894 9854 622338
rect 9234 586658 9266 586894
rect 9502 586658 9586 586894
rect 9822 586658 9854 586894
rect 9234 586574 9854 586658
rect 9234 586338 9266 586574
rect 9502 586338 9586 586574
rect 9822 586338 9854 586574
rect 9234 550894 9854 586338
rect 9234 550658 9266 550894
rect 9502 550658 9586 550894
rect 9822 550658 9854 550894
rect 9234 550574 9854 550658
rect 9234 550338 9266 550574
rect 9502 550338 9586 550574
rect 9822 550338 9854 550574
rect 9234 514894 9854 550338
rect 9234 514658 9266 514894
rect 9502 514658 9586 514894
rect 9822 514658 9854 514894
rect 9234 514574 9854 514658
rect 9234 514338 9266 514574
rect 9502 514338 9586 514574
rect 9822 514338 9854 514574
rect 9234 478894 9854 514338
rect 9234 478658 9266 478894
rect 9502 478658 9586 478894
rect 9822 478658 9854 478894
rect 9234 478574 9854 478658
rect 9234 478338 9266 478574
rect 9502 478338 9586 478574
rect 9822 478338 9854 478574
rect 9234 442894 9854 478338
rect 9234 442658 9266 442894
rect 9502 442658 9586 442894
rect 9822 442658 9854 442894
rect 9234 442574 9854 442658
rect 9234 442338 9266 442574
rect 9502 442338 9586 442574
rect 9822 442338 9854 442574
rect 9234 406894 9854 442338
rect 9234 406658 9266 406894
rect 9502 406658 9586 406894
rect 9822 406658 9854 406894
rect 9234 406574 9854 406658
rect 9234 406338 9266 406574
rect 9502 406338 9586 406574
rect 9822 406338 9854 406574
rect 9234 370894 9854 406338
rect 9234 370658 9266 370894
rect 9502 370658 9586 370894
rect 9822 370658 9854 370894
rect 9234 370574 9854 370658
rect 9234 370338 9266 370574
rect 9502 370338 9586 370574
rect 9822 370338 9854 370574
rect 9234 334894 9854 370338
rect 9234 334658 9266 334894
rect 9502 334658 9586 334894
rect 9822 334658 9854 334894
rect 9234 334574 9854 334658
rect 9234 334338 9266 334574
rect 9502 334338 9586 334574
rect 9822 334338 9854 334574
rect 9234 298894 9854 334338
rect 9234 298658 9266 298894
rect 9502 298658 9586 298894
rect 9822 298658 9854 298894
rect 9234 298574 9854 298658
rect 9234 298338 9266 298574
rect 9502 298338 9586 298574
rect 9822 298338 9854 298574
rect 9234 262894 9854 298338
rect 9234 262658 9266 262894
rect 9502 262658 9586 262894
rect 9822 262658 9854 262894
rect 9234 262574 9854 262658
rect 9234 262338 9266 262574
rect 9502 262338 9586 262574
rect 9822 262338 9854 262574
rect 9234 226894 9854 262338
rect 9234 226658 9266 226894
rect 9502 226658 9586 226894
rect 9822 226658 9854 226894
rect 9234 226574 9854 226658
rect 9234 226338 9266 226574
rect 9502 226338 9586 226574
rect 9822 226338 9854 226574
rect 9234 190894 9854 226338
rect 9234 190658 9266 190894
rect 9502 190658 9586 190894
rect 9822 190658 9854 190894
rect 9234 190574 9854 190658
rect 9234 190338 9266 190574
rect 9502 190338 9586 190574
rect 9822 190338 9854 190574
rect 9234 154894 9854 190338
rect 9234 154658 9266 154894
rect 9502 154658 9586 154894
rect 9822 154658 9854 154894
rect 9234 154574 9854 154658
rect 9234 154338 9266 154574
rect 9502 154338 9586 154574
rect 9822 154338 9854 154574
rect 9234 118894 9854 154338
rect 9234 118658 9266 118894
rect 9502 118658 9586 118894
rect 9822 118658 9854 118894
rect 9234 118574 9854 118658
rect 9234 118338 9266 118574
rect 9502 118338 9586 118574
rect 9822 118338 9854 118574
rect 9234 82894 9854 118338
rect 9234 82658 9266 82894
rect 9502 82658 9586 82894
rect 9822 82658 9854 82894
rect 9234 82574 9854 82658
rect 9234 82338 9266 82574
rect 9502 82338 9586 82574
rect 9822 82338 9854 82574
rect 9234 46894 9854 82338
rect 9234 46658 9266 46894
rect 9502 46658 9586 46894
rect 9822 46658 9854 46894
rect 9234 46574 9854 46658
rect 9234 46338 9266 46574
rect 9502 46338 9586 46574
rect 9822 46338 9854 46574
rect 9234 10894 9854 46338
rect 9234 10658 9266 10894
rect 9502 10658 9586 10894
rect 9822 10658 9854 10894
rect 9234 10574 9854 10658
rect 9234 10338 9266 10574
rect 9502 10338 9586 10574
rect 9822 10338 9854 10574
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 -5226 -4186
rect -5846 -4506 -5226 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 -5226 -4506
rect -5846 -4774 -5226 -4742
rect 9234 -4186 9854 10338
rect 9234 -4422 9266 -4186
rect 9502 -4422 9586 -4186
rect 9822 -4422 9854 -4186
rect 9234 -4506 9854 -4422
rect 9234 -4742 9266 -4506
rect 9502 -4742 9586 -4506
rect 9822 -4742 9854 -4506
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 -6186 -5146
rect -6806 -5466 -6186 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 -6186 -5466
rect -6806 -5734 -6186 -5702
rect 9234 -5734 9854 -4742
rect 12954 698614 13574 710042
rect 30954 711558 31574 711590
rect 30954 711322 30986 711558
rect 31222 711322 31306 711558
rect 31542 711322 31574 711558
rect 30954 711238 31574 711322
rect 30954 711002 30986 711238
rect 31222 711002 31306 711238
rect 31542 711002 31574 711238
rect 27234 709638 27854 709670
rect 27234 709402 27266 709638
rect 27502 709402 27586 709638
rect 27822 709402 27854 709638
rect 27234 709318 27854 709402
rect 27234 709082 27266 709318
rect 27502 709082 27586 709318
rect 27822 709082 27854 709318
rect 23514 707718 24134 707750
rect 23514 707482 23546 707718
rect 23782 707482 23866 707718
rect 24102 707482 24134 707718
rect 23514 707398 24134 707482
rect 23514 707162 23546 707398
rect 23782 707162 23866 707398
rect 24102 707162 24134 707398
rect 12954 698378 12986 698614
rect 13222 698378 13306 698614
rect 13542 698378 13574 698614
rect 12954 698294 13574 698378
rect 12954 698058 12986 698294
rect 13222 698058 13306 698294
rect 13542 698058 13574 698294
rect 12954 662614 13574 698058
rect 12954 662378 12986 662614
rect 13222 662378 13306 662614
rect 13542 662378 13574 662614
rect 12954 662294 13574 662378
rect 12954 662058 12986 662294
rect 13222 662058 13306 662294
rect 13542 662058 13574 662294
rect 12954 626614 13574 662058
rect 12954 626378 12986 626614
rect 13222 626378 13306 626614
rect 13542 626378 13574 626614
rect 12954 626294 13574 626378
rect 12954 626058 12986 626294
rect 13222 626058 13306 626294
rect 13542 626058 13574 626294
rect 12954 590614 13574 626058
rect 12954 590378 12986 590614
rect 13222 590378 13306 590614
rect 13542 590378 13574 590614
rect 12954 590294 13574 590378
rect 12954 590058 12986 590294
rect 13222 590058 13306 590294
rect 13542 590058 13574 590294
rect 12954 554614 13574 590058
rect 12954 554378 12986 554614
rect 13222 554378 13306 554614
rect 13542 554378 13574 554614
rect 12954 554294 13574 554378
rect 12954 554058 12986 554294
rect 13222 554058 13306 554294
rect 13542 554058 13574 554294
rect 12954 518614 13574 554058
rect 12954 518378 12986 518614
rect 13222 518378 13306 518614
rect 13542 518378 13574 518614
rect 12954 518294 13574 518378
rect 12954 518058 12986 518294
rect 13222 518058 13306 518294
rect 13542 518058 13574 518294
rect 12954 482614 13574 518058
rect 12954 482378 12986 482614
rect 13222 482378 13306 482614
rect 13542 482378 13574 482614
rect 12954 482294 13574 482378
rect 12954 482058 12986 482294
rect 13222 482058 13306 482294
rect 13542 482058 13574 482294
rect 12954 446614 13574 482058
rect 12954 446378 12986 446614
rect 13222 446378 13306 446614
rect 13542 446378 13574 446614
rect 12954 446294 13574 446378
rect 12954 446058 12986 446294
rect 13222 446058 13306 446294
rect 13542 446058 13574 446294
rect 12954 410614 13574 446058
rect 12954 410378 12986 410614
rect 13222 410378 13306 410614
rect 13542 410378 13574 410614
rect 12954 410294 13574 410378
rect 12954 410058 12986 410294
rect 13222 410058 13306 410294
rect 13542 410058 13574 410294
rect 12954 374614 13574 410058
rect 12954 374378 12986 374614
rect 13222 374378 13306 374614
rect 13542 374378 13574 374614
rect 12954 374294 13574 374378
rect 12954 374058 12986 374294
rect 13222 374058 13306 374294
rect 13542 374058 13574 374294
rect 12954 338614 13574 374058
rect 12954 338378 12986 338614
rect 13222 338378 13306 338614
rect 13542 338378 13574 338614
rect 12954 338294 13574 338378
rect 12954 338058 12986 338294
rect 13222 338058 13306 338294
rect 13542 338058 13574 338294
rect 12954 302614 13574 338058
rect 12954 302378 12986 302614
rect 13222 302378 13306 302614
rect 13542 302378 13574 302614
rect 12954 302294 13574 302378
rect 12954 302058 12986 302294
rect 13222 302058 13306 302294
rect 13542 302058 13574 302294
rect 12954 266614 13574 302058
rect 12954 266378 12986 266614
rect 13222 266378 13306 266614
rect 13542 266378 13574 266614
rect 12954 266294 13574 266378
rect 12954 266058 12986 266294
rect 13222 266058 13306 266294
rect 13542 266058 13574 266294
rect 12954 230614 13574 266058
rect 12954 230378 12986 230614
rect 13222 230378 13306 230614
rect 13542 230378 13574 230614
rect 12954 230294 13574 230378
rect 12954 230058 12986 230294
rect 13222 230058 13306 230294
rect 13542 230058 13574 230294
rect 12954 194614 13574 230058
rect 12954 194378 12986 194614
rect 13222 194378 13306 194614
rect 13542 194378 13574 194614
rect 12954 194294 13574 194378
rect 12954 194058 12986 194294
rect 13222 194058 13306 194294
rect 13542 194058 13574 194294
rect 12954 158614 13574 194058
rect 12954 158378 12986 158614
rect 13222 158378 13306 158614
rect 13542 158378 13574 158614
rect 12954 158294 13574 158378
rect 12954 158058 12986 158294
rect 13222 158058 13306 158294
rect 13542 158058 13574 158294
rect 12954 122614 13574 158058
rect 12954 122378 12986 122614
rect 13222 122378 13306 122614
rect 13542 122378 13574 122614
rect 12954 122294 13574 122378
rect 12954 122058 12986 122294
rect 13222 122058 13306 122294
rect 13542 122058 13574 122294
rect 12954 86614 13574 122058
rect 12954 86378 12986 86614
rect 13222 86378 13306 86614
rect 13542 86378 13574 86614
rect 12954 86294 13574 86378
rect 12954 86058 12986 86294
rect 13222 86058 13306 86294
rect 13542 86058 13574 86294
rect 12954 50614 13574 86058
rect 12954 50378 12986 50614
rect 13222 50378 13306 50614
rect 13542 50378 13574 50614
rect 12954 50294 13574 50378
rect 12954 50058 12986 50294
rect 13222 50058 13306 50294
rect 13542 50058 13574 50294
rect 12954 14614 13574 50058
rect 12954 14378 12986 14614
rect 13222 14378 13306 14614
rect 13542 14378 13574 14614
rect 12954 14294 13574 14378
rect 12954 14058 12986 14294
rect 13222 14058 13306 14294
rect 13542 14058 13574 14294
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 -7146 -6106
rect -7766 -6426 -7146 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 -7146 -6426
rect -7766 -6694 -7146 -6662
rect 12954 -6106 13574 14058
rect 19794 705798 20414 705830
rect 19794 705562 19826 705798
rect 20062 705562 20146 705798
rect 20382 705562 20414 705798
rect 19794 705478 20414 705562
rect 19794 705242 19826 705478
rect 20062 705242 20146 705478
rect 20382 705242 20414 705478
rect 19794 669454 20414 705242
rect 19794 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 20414 669454
rect 19794 669134 20414 669218
rect 19794 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 20414 669134
rect 19794 633454 20414 668898
rect 19794 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 20414 633454
rect 19794 633134 20414 633218
rect 19794 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 20414 633134
rect 19794 597454 20414 632898
rect 19794 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 20414 597454
rect 19794 597134 20414 597218
rect 19794 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 20414 597134
rect 19794 561454 20414 596898
rect 19794 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 20414 561454
rect 19794 561134 20414 561218
rect 19794 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 20414 561134
rect 19794 525454 20414 560898
rect 19794 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 20414 525454
rect 19794 525134 20414 525218
rect 19794 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 20414 525134
rect 19794 489454 20414 524898
rect 19794 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 20414 489454
rect 19794 489134 20414 489218
rect 19794 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 20414 489134
rect 19794 453454 20414 488898
rect 19794 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 20414 453454
rect 19794 453134 20414 453218
rect 19794 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 20414 453134
rect 19794 417454 20414 452898
rect 19794 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 20414 417454
rect 19794 417134 20414 417218
rect 19794 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 20414 417134
rect 19794 381454 20414 416898
rect 19794 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 20414 381454
rect 19794 381134 20414 381218
rect 19794 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 20414 381134
rect 19794 345454 20414 380898
rect 19794 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 20414 345454
rect 19794 345134 20414 345218
rect 19794 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 20414 345134
rect 19794 309454 20414 344898
rect 19794 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 20414 309454
rect 19794 309134 20414 309218
rect 19794 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 20414 309134
rect 19794 273454 20414 308898
rect 19794 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 20414 273454
rect 19794 273134 20414 273218
rect 19794 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 20414 273134
rect 19794 237454 20414 272898
rect 19794 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 20414 237454
rect 19794 237134 20414 237218
rect 19794 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 20414 237134
rect 19794 201454 20414 236898
rect 19794 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 20414 201454
rect 19794 201134 20414 201218
rect 19794 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 20414 201134
rect 19794 165454 20414 200898
rect 19794 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 20414 165454
rect 19794 165134 20414 165218
rect 19794 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 20414 165134
rect 19794 129454 20414 164898
rect 19794 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 20414 129454
rect 19794 129134 20414 129218
rect 19794 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 20414 129134
rect 19794 93454 20414 128898
rect 19794 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 20414 93454
rect 19794 93134 20414 93218
rect 19794 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 20414 93134
rect 19794 57454 20414 92898
rect 19794 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 20414 57454
rect 19794 57134 20414 57218
rect 19794 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 20414 57134
rect 19794 21454 20414 56898
rect 19794 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 20414 21454
rect 19794 21134 20414 21218
rect 19794 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 20414 21134
rect 19794 -1306 20414 20898
rect 19794 -1542 19826 -1306
rect 20062 -1542 20146 -1306
rect 20382 -1542 20414 -1306
rect 19794 -1626 20414 -1542
rect 19794 -1862 19826 -1626
rect 20062 -1862 20146 -1626
rect 20382 -1862 20414 -1626
rect 19794 -1894 20414 -1862
rect 23514 673174 24134 707162
rect 23514 672938 23546 673174
rect 23782 672938 23866 673174
rect 24102 672938 24134 673174
rect 23514 672854 24134 672938
rect 23514 672618 23546 672854
rect 23782 672618 23866 672854
rect 24102 672618 24134 672854
rect 23514 637174 24134 672618
rect 23514 636938 23546 637174
rect 23782 636938 23866 637174
rect 24102 636938 24134 637174
rect 23514 636854 24134 636938
rect 23514 636618 23546 636854
rect 23782 636618 23866 636854
rect 24102 636618 24134 636854
rect 23514 601174 24134 636618
rect 23514 600938 23546 601174
rect 23782 600938 23866 601174
rect 24102 600938 24134 601174
rect 23514 600854 24134 600938
rect 23514 600618 23546 600854
rect 23782 600618 23866 600854
rect 24102 600618 24134 600854
rect 23514 565174 24134 600618
rect 23514 564938 23546 565174
rect 23782 564938 23866 565174
rect 24102 564938 24134 565174
rect 23514 564854 24134 564938
rect 23514 564618 23546 564854
rect 23782 564618 23866 564854
rect 24102 564618 24134 564854
rect 23514 529174 24134 564618
rect 23514 528938 23546 529174
rect 23782 528938 23866 529174
rect 24102 528938 24134 529174
rect 23514 528854 24134 528938
rect 23514 528618 23546 528854
rect 23782 528618 23866 528854
rect 24102 528618 24134 528854
rect 23514 493174 24134 528618
rect 23514 492938 23546 493174
rect 23782 492938 23866 493174
rect 24102 492938 24134 493174
rect 23514 492854 24134 492938
rect 23514 492618 23546 492854
rect 23782 492618 23866 492854
rect 24102 492618 24134 492854
rect 23514 457174 24134 492618
rect 23514 456938 23546 457174
rect 23782 456938 23866 457174
rect 24102 456938 24134 457174
rect 23514 456854 24134 456938
rect 23514 456618 23546 456854
rect 23782 456618 23866 456854
rect 24102 456618 24134 456854
rect 23514 421174 24134 456618
rect 23514 420938 23546 421174
rect 23782 420938 23866 421174
rect 24102 420938 24134 421174
rect 23514 420854 24134 420938
rect 23514 420618 23546 420854
rect 23782 420618 23866 420854
rect 24102 420618 24134 420854
rect 23514 385174 24134 420618
rect 23514 384938 23546 385174
rect 23782 384938 23866 385174
rect 24102 384938 24134 385174
rect 23514 384854 24134 384938
rect 23514 384618 23546 384854
rect 23782 384618 23866 384854
rect 24102 384618 24134 384854
rect 23514 349174 24134 384618
rect 23514 348938 23546 349174
rect 23782 348938 23866 349174
rect 24102 348938 24134 349174
rect 23514 348854 24134 348938
rect 23514 348618 23546 348854
rect 23782 348618 23866 348854
rect 24102 348618 24134 348854
rect 23514 313174 24134 348618
rect 23514 312938 23546 313174
rect 23782 312938 23866 313174
rect 24102 312938 24134 313174
rect 23514 312854 24134 312938
rect 23514 312618 23546 312854
rect 23782 312618 23866 312854
rect 24102 312618 24134 312854
rect 23514 277174 24134 312618
rect 23514 276938 23546 277174
rect 23782 276938 23866 277174
rect 24102 276938 24134 277174
rect 23514 276854 24134 276938
rect 23514 276618 23546 276854
rect 23782 276618 23866 276854
rect 24102 276618 24134 276854
rect 23514 241174 24134 276618
rect 23514 240938 23546 241174
rect 23782 240938 23866 241174
rect 24102 240938 24134 241174
rect 23514 240854 24134 240938
rect 23514 240618 23546 240854
rect 23782 240618 23866 240854
rect 24102 240618 24134 240854
rect 23514 205174 24134 240618
rect 23514 204938 23546 205174
rect 23782 204938 23866 205174
rect 24102 204938 24134 205174
rect 23514 204854 24134 204938
rect 23514 204618 23546 204854
rect 23782 204618 23866 204854
rect 24102 204618 24134 204854
rect 23514 169174 24134 204618
rect 23514 168938 23546 169174
rect 23782 168938 23866 169174
rect 24102 168938 24134 169174
rect 23514 168854 24134 168938
rect 23514 168618 23546 168854
rect 23782 168618 23866 168854
rect 24102 168618 24134 168854
rect 23514 133174 24134 168618
rect 23514 132938 23546 133174
rect 23782 132938 23866 133174
rect 24102 132938 24134 133174
rect 23514 132854 24134 132938
rect 23514 132618 23546 132854
rect 23782 132618 23866 132854
rect 24102 132618 24134 132854
rect 23514 97174 24134 132618
rect 23514 96938 23546 97174
rect 23782 96938 23866 97174
rect 24102 96938 24134 97174
rect 23514 96854 24134 96938
rect 23514 96618 23546 96854
rect 23782 96618 23866 96854
rect 24102 96618 24134 96854
rect 23514 61174 24134 96618
rect 23514 60938 23546 61174
rect 23782 60938 23866 61174
rect 24102 60938 24134 61174
rect 23514 60854 24134 60938
rect 23514 60618 23546 60854
rect 23782 60618 23866 60854
rect 24102 60618 24134 60854
rect 23514 25174 24134 60618
rect 23514 24938 23546 25174
rect 23782 24938 23866 25174
rect 24102 24938 24134 25174
rect 23514 24854 24134 24938
rect 23514 24618 23546 24854
rect 23782 24618 23866 24854
rect 24102 24618 24134 24854
rect 23514 -3226 24134 24618
rect 23514 -3462 23546 -3226
rect 23782 -3462 23866 -3226
rect 24102 -3462 24134 -3226
rect 23514 -3546 24134 -3462
rect 23514 -3782 23546 -3546
rect 23782 -3782 23866 -3546
rect 24102 -3782 24134 -3546
rect 23514 -3814 24134 -3782
rect 27234 676894 27854 709082
rect 27234 676658 27266 676894
rect 27502 676658 27586 676894
rect 27822 676658 27854 676894
rect 27234 676574 27854 676658
rect 27234 676338 27266 676574
rect 27502 676338 27586 676574
rect 27822 676338 27854 676574
rect 27234 640894 27854 676338
rect 27234 640658 27266 640894
rect 27502 640658 27586 640894
rect 27822 640658 27854 640894
rect 27234 640574 27854 640658
rect 27234 640338 27266 640574
rect 27502 640338 27586 640574
rect 27822 640338 27854 640574
rect 27234 604894 27854 640338
rect 27234 604658 27266 604894
rect 27502 604658 27586 604894
rect 27822 604658 27854 604894
rect 27234 604574 27854 604658
rect 27234 604338 27266 604574
rect 27502 604338 27586 604574
rect 27822 604338 27854 604574
rect 27234 568894 27854 604338
rect 27234 568658 27266 568894
rect 27502 568658 27586 568894
rect 27822 568658 27854 568894
rect 27234 568574 27854 568658
rect 27234 568338 27266 568574
rect 27502 568338 27586 568574
rect 27822 568338 27854 568574
rect 27234 532894 27854 568338
rect 27234 532658 27266 532894
rect 27502 532658 27586 532894
rect 27822 532658 27854 532894
rect 27234 532574 27854 532658
rect 27234 532338 27266 532574
rect 27502 532338 27586 532574
rect 27822 532338 27854 532574
rect 27234 496894 27854 532338
rect 27234 496658 27266 496894
rect 27502 496658 27586 496894
rect 27822 496658 27854 496894
rect 27234 496574 27854 496658
rect 27234 496338 27266 496574
rect 27502 496338 27586 496574
rect 27822 496338 27854 496574
rect 27234 460894 27854 496338
rect 27234 460658 27266 460894
rect 27502 460658 27586 460894
rect 27822 460658 27854 460894
rect 27234 460574 27854 460658
rect 27234 460338 27266 460574
rect 27502 460338 27586 460574
rect 27822 460338 27854 460574
rect 27234 424894 27854 460338
rect 27234 424658 27266 424894
rect 27502 424658 27586 424894
rect 27822 424658 27854 424894
rect 27234 424574 27854 424658
rect 27234 424338 27266 424574
rect 27502 424338 27586 424574
rect 27822 424338 27854 424574
rect 27234 388894 27854 424338
rect 27234 388658 27266 388894
rect 27502 388658 27586 388894
rect 27822 388658 27854 388894
rect 27234 388574 27854 388658
rect 27234 388338 27266 388574
rect 27502 388338 27586 388574
rect 27822 388338 27854 388574
rect 27234 352894 27854 388338
rect 27234 352658 27266 352894
rect 27502 352658 27586 352894
rect 27822 352658 27854 352894
rect 27234 352574 27854 352658
rect 27234 352338 27266 352574
rect 27502 352338 27586 352574
rect 27822 352338 27854 352574
rect 27234 316894 27854 352338
rect 27234 316658 27266 316894
rect 27502 316658 27586 316894
rect 27822 316658 27854 316894
rect 27234 316574 27854 316658
rect 27234 316338 27266 316574
rect 27502 316338 27586 316574
rect 27822 316338 27854 316574
rect 27234 280894 27854 316338
rect 27234 280658 27266 280894
rect 27502 280658 27586 280894
rect 27822 280658 27854 280894
rect 27234 280574 27854 280658
rect 27234 280338 27266 280574
rect 27502 280338 27586 280574
rect 27822 280338 27854 280574
rect 27234 244894 27854 280338
rect 27234 244658 27266 244894
rect 27502 244658 27586 244894
rect 27822 244658 27854 244894
rect 27234 244574 27854 244658
rect 27234 244338 27266 244574
rect 27502 244338 27586 244574
rect 27822 244338 27854 244574
rect 27234 208894 27854 244338
rect 27234 208658 27266 208894
rect 27502 208658 27586 208894
rect 27822 208658 27854 208894
rect 27234 208574 27854 208658
rect 27234 208338 27266 208574
rect 27502 208338 27586 208574
rect 27822 208338 27854 208574
rect 27234 172894 27854 208338
rect 27234 172658 27266 172894
rect 27502 172658 27586 172894
rect 27822 172658 27854 172894
rect 27234 172574 27854 172658
rect 27234 172338 27266 172574
rect 27502 172338 27586 172574
rect 27822 172338 27854 172574
rect 27234 136894 27854 172338
rect 27234 136658 27266 136894
rect 27502 136658 27586 136894
rect 27822 136658 27854 136894
rect 27234 136574 27854 136658
rect 27234 136338 27266 136574
rect 27502 136338 27586 136574
rect 27822 136338 27854 136574
rect 27234 100894 27854 136338
rect 27234 100658 27266 100894
rect 27502 100658 27586 100894
rect 27822 100658 27854 100894
rect 27234 100574 27854 100658
rect 27234 100338 27266 100574
rect 27502 100338 27586 100574
rect 27822 100338 27854 100574
rect 27234 64894 27854 100338
rect 27234 64658 27266 64894
rect 27502 64658 27586 64894
rect 27822 64658 27854 64894
rect 27234 64574 27854 64658
rect 27234 64338 27266 64574
rect 27502 64338 27586 64574
rect 27822 64338 27854 64574
rect 27234 28894 27854 64338
rect 27234 28658 27266 28894
rect 27502 28658 27586 28894
rect 27822 28658 27854 28894
rect 27234 28574 27854 28658
rect 27234 28338 27266 28574
rect 27502 28338 27586 28574
rect 27822 28338 27854 28574
rect 27234 -5146 27854 28338
rect 27234 -5382 27266 -5146
rect 27502 -5382 27586 -5146
rect 27822 -5382 27854 -5146
rect 27234 -5466 27854 -5382
rect 27234 -5702 27266 -5466
rect 27502 -5702 27586 -5466
rect 27822 -5702 27854 -5466
rect 27234 -5734 27854 -5702
rect 30954 680614 31574 711002
rect 48954 710598 49574 711590
rect 48954 710362 48986 710598
rect 49222 710362 49306 710598
rect 49542 710362 49574 710598
rect 48954 710278 49574 710362
rect 48954 710042 48986 710278
rect 49222 710042 49306 710278
rect 49542 710042 49574 710278
rect 45234 708678 45854 709670
rect 45234 708442 45266 708678
rect 45502 708442 45586 708678
rect 45822 708442 45854 708678
rect 45234 708358 45854 708442
rect 45234 708122 45266 708358
rect 45502 708122 45586 708358
rect 45822 708122 45854 708358
rect 41514 706758 42134 707750
rect 41514 706522 41546 706758
rect 41782 706522 41866 706758
rect 42102 706522 42134 706758
rect 41514 706438 42134 706522
rect 41514 706202 41546 706438
rect 41782 706202 41866 706438
rect 42102 706202 42134 706438
rect 30954 680378 30986 680614
rect 31222 680378 31306 680614
rect 31542 680378 31574 680614
rect 30954 680294 31574 680378
rect 30954 680058 30986 680294
rect 31222 680058 31306 680294
rect 31542 680058 31574 680294
rect 30954 644614 31574 680058
rect 30954 644378 30986 644614
rect 31222 644378 31306 644614
rect 31542 644378 31574 644614
rect 30954 644294 31574 644378
rect 30954 644058 30986 644294
rect 31222 644058 31306 644294
rect 31542 644058 31574 644294
rect 30954 608614 31574 644058
rect 30954 608378 30986 608614
rect 31222 608378 31306 608614
rect 31542 608378 31574 608614
rect 30954 608294 31574 608378
rect 30954 608058 30986 608294
rect 31222 608058 31306 608294
rect 31542 608058 31574 608294
rect 30954 572614 31574 608058
rect 30954 572378 30986 572614
rect 31222 572378 31306 572614
rect 31542 572378 31574 572614
rect 30954 572294 31574 572378
rect 30954 572058 30986 572294
rect 31222 572058 31306 572294
rect 31542 572058 31574 572294
rect 30954 536614 31574 572058
rect 30954 536378 30986 536614
rect 31222 536378 31306 536614
rect 31542 536378 31574 536614
rect 30954 536294 31574 536378
rect 30954 536058 30986 536294
rect 31222 536058 31306 536294
rect 31542 536058 31574 536294
rect 30954 500614 31574 536058
rect 30954 500378 30986 500614
rect 31222 500378 31306 500614
rect 31542 500378 31574 500614
rect 30954 500294 31574 500378
rect 30954 500058 30986 500294
rect 31222 500058 31306 500294
rect 31542 500058 31574 500294
rect 30954 464614 31574 500058
rect 30954 464378 30986 464614
rect 31222 464378 31306 464614
rect 31542 464378 31574 464614
rect 30954 464294 31574 464378
rect 30954 464058 30986 464294
rect 31222 464058 31306 464294
rect 31542 464058 31574 464294
rect 30954 428614 31574 464058
rect 30954 428378 30986 428614
rect 31222 428378 31306 428614
rect 31542 428378 31574 428614
rect 30954 428294 31574 428378
rect 30954 428058 30986 428294
rect 31222 428058 31306 428294
rect 31542 428058 31574 428294
rect 30954 392614 31574 428058
rect 30954 392378 30986 392614
rect 31222 392378 31306 392614
rect 31542 392378 31574 392614
rect 30954 392294 31574 392378
rect 30954 392058 30986 392294
rect 31222 392058 31306 392294
rect 31542 392058 31574 392294
rect 30954 356614 31574 392058
rect 30954 356378 30986 356614
rect 31222 356378 31306 356614
rect 31542 356378 31574 356614
rect 30954 356294 31574 356378
rect 30954 356058 30986 356294
rect 31222 356058 31306 356294
rect 31542 356058 31574 356294
rect 30954 320614 31574 356058
rect 30954 320378 30986 320614
rect 31222 320378 31306 320614
rect 31542 320378 31574 320614
rect 30954 320294 31574 320378
rect 30954 320058 30986 320294
rect 31222 320058 31306 320294
rect 31542 320058 31574 320294
rect 30954 284614 31574 320058
rect 30954 284378 30986 284614
rect 31222 284378 31306 284614
rect 31542 284378 31574 284614
rect 30954 284294 31574 284378
rect 30954 284058 30986 284294
rect 31222 284058 31306 284294
rect 31542 284058 31574 284294
rect 30954 248614 31574 284058
rect 30954 248378 30986 248614
rect 31222 248378 31306 248614
rect 31542 248378 31574 248614
rect 30954 248294 31574 248378
rect 30954 248058 30986 248294
rect 31222 248058 31306 248294
rect 31542 248058 31574 248294
rect 30954 212614 31574 248058
rect 30954 212378 30986 212614
rect 31222 212378 31306 212614
rect 31542 212378 31574 212614
rect 30954 212294 31574 212378
rect 30954 212058 30986 212294
rect 31222 212058 31306 212294
rect 31542 212058 31574 212294
rect 30954 176614 31574 212058
rect 30954 176378 30986 176614
rect 31222 176378 31306 176614
rect 31542 176378 31574 176614
rect 30954 176294 31574 176378
rect 30954 176058 30986 176294
rect 31222 176058 31306 176294
rect 31542 176058 31574 176294
rect 30954 140614 31574 176058
rect 30954 140378 30986 140614
rect 31222 140378 31306 140614
rect 31542 140378 31574 140614
rect 30954 140294 31574 140378
rect 30954 140058 30986 140294
rect 31222 140058 31306 140294
rect 31542 140058 31574 140294
rect 30954 104614 31574 140058
rect 30954 104378 30986 104614
rect 31222 104378 31306 104614
rect 31542 104378 31574 104614
rect 30954 104294 31574 104378
rect 30954 104058 30986 104294
rect 31222 104058 31306 104294
rect 31542 104058 31574 104294
rect 30954 68614 31574 104058
rect 30954 68378 30986 68614
rect 31222 68378 31306 68614
rect 31542 68378 31574 68614
rect 30954 68294 31574 68378
rect 30954 68058 30986 68294
rect 31222 68058 31306 68294
rect 31542 68058 31574 68294
rect 30954 32614 31574 68058
rect 30954 32378 30986 32614
rect 31222 32378 31306 32614
rect 31542 32378 31574 32614
rect 30954 32294 31574 32378
rect 30954 32058 30986 32294
rect 31222 32058 31306 32294
rect 31542 32058 31574 32294
rect 12954 -6342 12986 -6106
rect 13222 -6342 13306 -6106
rect 13542 -6342 13574 -6106
rect 12954 -6426 13574 -6342
rect 12954 -6662 12986 -6426
rect 13222 -6662 13306 -6426
rect 13542 -6662 13574 -6426
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 -8106 -7066
rect -8726 -7386 -8106 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 -8106 -7386
rect -8726 -7654 -8106 -7622
rect 12954 -7654 13574 -6662
rect 30954 -7066 31574 32058
rect 37794 704838 38414 705830
rect 37794 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 38414 704838
rect 37794 704518 38414 704602
rect 37794 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 38414 704518
rect 37794 687454 38414 704282
rect 37794 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 38414 687454
rect 37794 687134 38414 687218
rect 37794 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 38414 687134
rect 37794 651454 38414 686898
rect 37794 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 38414 651454
rect 37794 651134 38414 651218
rect 37794 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 38414 651134
rect 37794 615454 38414 650898
rect 37794 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 38414 615454
rect 37794 615134 38414 615218
rect 37794 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 38414 615134
rect 37794 579454 38414 614898
rect 37794 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 38414 579454
rect 37794 579134 38414 579218
rect 37794 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 38414 579134
rect 37794 543454 38414 578898
rect 37794 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 38414 543454
rect 37794 543134 38414 543218
rect 37794 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 38414 543134
rect 37794 507454 38414 542898
rect 37794 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 38414 507454
rect 37794 507134 38414 507218
rect 37794 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 38414 507134
rect 37794 471454 38414 506898
rect 37794 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 38414 471454
rect 37794 471134 38414 471218
rect 37794 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 38414 471134
rect 37794 435454 38414 470898
rect 37794 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 38414 435454
rect 37794 435134 38414 435218
rect 37794 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 38414 435134
rect 37794 399454 38414 434898
rect 37794 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 38414 399454
rect 37794 399134 38414 399218
rect 37794 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 38414 399134
rect 37794 363454 38414 398898
rect 37794 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 38414 363454
rect 37794 363134 38414 363218
rect 37794 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 38414 363134
rect 37794 327454 38414 362898
rect 37794 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 38414 327454
rect 37794 327134 38414 327218
rect 37794 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 38414 327134
rect 37794 291454 38414 326898
rect 37794 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 38414 291454
rect 37794 291134 38414 291218
rect 37794 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 38414 291134
rect 37794 255454 38414 290898
rect 37794 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 38414 255454
rect 37794 255134 38414 255218
rect 37794 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 38414 255134
rect 37794 219454 38414 254898
rect 37794 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 38414 219454
rect 37794 219134 38414 219218
rect 37794 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 38414 219134
rect 37794 183454 38414 218898
rect 37794 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 38414 183454
rect 37794 183134 38414 183218
rect 37794 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 38414 183134
rect 37794 147454 38414 182898
rect 37794 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 38414 147454
rect 37794 147134 38414 147218
rect 37794 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 38414 147134
rect 37794 111454 38414 146898
rect 37794 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 38414 111454
rect 37794 111134 38414 111218
rect 37794 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 38414 111134
rect 37794 75454 38414 110898
rect 37794 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 38414 75454
rect 37794 75134 38414 75218
rect 37794 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 38414 75134
rect 37794 39454 38414 74898
rect 37794 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 38414 39454
rect 37794 39134 38414 39218
rect 37794 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 38414 39134
rect 37794 3454 38414 38898
rect 37794 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 38414 3454
rect 37794 3134 38414 3218
rect 37794 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 38414 3134
rect 37794 -346 38414 2898
rect 37794 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 38414 -346
rect 37794 -666 38414 -582
rect 37794 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 38414 -666
rect 37794 -1894 38414 -902
rect 41514 691174 42134 706202
rect 41514 690938 41546 691174
rect 41782 690938 41866 691174
rect 42102 690938 42134 691174
rect 41514 690854 42134 690938
rect 41514 690618 41546 690854
rect 41782 690618 41866 690854
rect 42102 690618 42134 690854
rect 41514 655174 42134 690618
rect 41514 654938 41546 655174
rect 41782 654938 41866 655174
rect 42102 654938 42134 655174
rect 41514 654854 42134 654938
rect 41514 654618 41546 654854
rect 41782 654618 41866 654854
rect 42102 654618 42134 654854
rect 41514 619174 42134 654618
rect 41514 618938 41546 619174
rect 41782 618938 41866 619174
rect 42102 618938 42134 619174
rect 41514 618854 42134 618938
rect 41514 618618 41546 618854
rect 41782 618618 41866 618854
rect 42102 618618 42134 618854
rect 41514 583174 42134 618618
rect 41514 582938 41546 583174
rect 41782 582938 41866 583174
rect 42102 582938 42134 583174
rect 41514 582854 42134 582938
rect 41514 582618 41546 582854
rect 41782 582618 41866 582854
rect 42102 582618 42134 582854
rect 41514 547174 42134 582618
rect 41514 546938 41546 547174
rect 41782 546938 41866 547174
rect 42102 546938 42134 547174
rect 41514 546854 42134 546938
rect 41514 546618 41546 546854
rect 41782 546618 41866 546854
rect 42102 546618 42134 546854
rect 41514 511174 42134 546618
rect 41514 510938 41546 511174
rect 41782 510938 41866 511174
rect 42102 510938 42134 511174
rect 41514 510854 42134 510938
rect 41514 510618 41546 510854
rect 41782 510618 41866 510854
rect 42102 510618 42134 510854
rect 41514 475174 42134 510618
rect 41514 474938 41546 475174
rect 41782 474938 41866 475174
rect 42102 474938 42134 475174
rect 41514 474854 42134 474938
rect 41514 474618 41546 474854
rect 41782 474618 41866 474854
rect 42102 474618 42134 474854
rect 41514 439174 42134 474618
rect 41514 438938 41546 439174
rect 41782 438938 41866 439174
rect 42102 438938 42134 439174
rect 41514 438854 42134 438938
rect 41514 438618 41546 438854
rect 41782 438618 41866 438854
rect 42102 438618 42134 438854
rect 41514 403174 42134 438618
rect 41514 402938 41546 403174
rect 41782 402938 41866 403174
rect 42102 402938 42134 403174
rect 41514 402854 42134 402938
rect 41514 402618 41546 402854
rect 41782 402618 41866 402854
rect 42102 402618 42134 402854
rect 41514 367174 42134 402618
rect 41514 366938 41546 367174
rect 41782 366938 41866 367174
rect 42102 366938 42134 367174
rect 41514 366854 42134 366938
rect 41514 366618 41546 366854
rect 41782 366618 41866 366854
rect 42102 366618 42134 366854
rect 41514 331174 42134 366618
rect 41514 330938 41546 331174
rect 41782 330938 41866 331174
rect 42102 330938 42134 331174
rect 41514 330854 42134 330938
rect 41514 330618 41546 330854
rect 41782 330618 41866 330854
rect 42102 330618 42134 330854
rect 41514 295174 42134 330618
rect 41514 294938 41546 295174
rect 41782 294938 41866 295174
rect 42102 294938 42134 295174
rect 41514 294854 42134 294938
rect 41514 294618 41546 294854
rect 41782 294618 41866 294854
rect 42102 294618 42134 294854
rect 41514 259174 42134 294618
rect 41514 258938 41546 259174
rect 41782 258938 41866 259174
rect 42102 258938 42134 259174
rect 41514 258854 42134 258938
rect 41514 258618 41546 258854
rect 41782 258618 41866 258854
rect 42102 258618 42134 258854
rect 41514 223174 42134 258618
rect 41514 222938 41546 223174
rect 41782 222938 41866 223174
rect 42102 222938 42134 223174
rect 41514 222854 42134 222938
rect 41514 222618 41546 222854
rect 41782 222618 41866 222854
rect 42102 222618 42134 222854
rect 41514 187174 42134 222618
rect 41514 186938 41546 187174
rect 41782 186938 41866 187174
rect 42102 186938 42134 187174
rect 41514 186854 42134 186938
rect 41514 186618 41546 186854
rect 41782 186618 41866 186854
rect 42102 186618 42134 186854
rect 41514 151174 42134 186618
rect 41514 150938 41546 151174
rect 41782 150938 41866 151174
rect 42102 150938 42134 151174
rect 41514 150854 42134 150938
rect 41514 150618 41546 150854
rect 41782 150618 41866 150854
rect 42102 150618 42134 150854
rect 41514 115174 42134 150618
rect 41514 114938 41546 115174
rect 41782 114938 41866 115174
rect 42102 114938 42134 115174
rect 41514 114854 42134 114938
rect 41514 114618 41546 114854
rect 41782 114618 41866 114854
rect 42102 114618 42134 114854
rect 41514 79174 42134 114618
rect 41514 78938 41546 79174
rect 41782 78938 41866 79174
rect 42102 78938 42134 79174
rect 41514 78854 42134 78938
rect 41514 78618 41546 78854
rect 41782 78618 41866 78854
rect 42102 78618 42134 78854
rect 41514 43174 42134 78618
rect 41514 42938 41546 43174
rect 41782 42938 41866 43174
rect 42102 42938 42134 43174
rect 41514 42854 42134 42938
rect 41514 42618 41546 42854
rect 41782 42618 41866 42854
rect 42102 42618 42134 42854
rect 41514 7174 42134 42618
rect 41514 6938 41546 7174
rect 41782 6938 41866 7174
rect 42102 6938 42134 7174
rect 41514 6854 42134 6938
rect 41514 6618 41546 6854
rect 41782 6618 41866 6854
rect 42102 6618 42134 6854
rect 41514 -2266 42134 6618
rect 41514 -2502 41546 -2266
rect 41782 -2502 41866 -2266
rect 42102 -2502 42134 -2266
rect 41514 -2586 42134 -2502
rect 41514 -2822 41546 -2586
rect 41782 -2822 41866 -2586
rect 42102 -2822 42134 -2586
rect 41514 -3814 42134 -2822
rect 45234 694894 45854 708122
rect 45234 694658 45266 694894
rect 45502 694658 45586 694894
rect 45822 694658 45854 694894
rect 45234 694574 45854 694658
rect 45234 694338 45266 694574
rect 45502 694338 45586 694574
rect 45822 694338 45854 694574
rect 45234 658894 45854 694338
rect 45234 658658 45266 658894
rect 45502 658658 45586 658894
rect 45822 658658 45854 658894
rect 45234 658574 45854 658658
rect 45234 658338 45266 658574
rect 45502 658338 45586 658574
rect 45822 658338 45854 658574
rect 45234 622894 45854 658338
rect 45234 622658 45266 622894
rect 45502 622658 45586 622894
rect 45822 622658 45854 622894
rect 45234 622574 45854 622658
rect 45234 622338 45266 622574
rect 45502 622338 45586 622574
rect 45822 622338 45854 622574
rect 45234 586894 45854 622338
rect 45234 586658 45266 586894
rect 45502 586658 45586 586894
rect 45822 586658 45854 586894
rect 45234 586574 45854 586658
rect 45234 586338 45266 586574
rect 45502 586338 45586 586574
rect 45822 586338 45854 586574
rect 45234 550894 45854 586338
rect 45234 550658 45266 550894
rect 45502 550658 45586 550894
rect 45822 550658 45854 550894
rect 45234 550574 45854 550658
rect 45234 550338 45266 550574
rect 45502 550338 45586 550574
rect 45822 550338 45854 550574
rect 45234 514894 45854 550338
rect 45234 514658 45266 514894
rect 45502 514658 45586 514894
rect 45822 514658 45854 514894
rect 45234 514574 45854 514658
rect 45234 514338 45266 514574
rect 45502 514338 45586 514574
rect 45822 514338 45854 514574
rect 45234 478894 45854 514338
rect 45234 478658 45266 478894
rect 45502 478658 45586 478894
rect 45822 478658 45854 478894
rect 45234 478574 45854 478658
rect 45234 478338 45266 478574
rect 45502 478338 45586 478574
rect 45822 478338 45854 478574
rect 45234 442894 45854 478338
rect 45234 442658 45266 442894
rect 45502 442658 45586 442894
rect 45822 442658 45854 442894
rect 45234 442574 45854 442658
rect 45234 442338 45266 442574
rect 45502 442338 45586 442574
rect 45822 442338 45854 442574
rect 45234 406894 45854 442338
rect 45234 406658 45266 406894
rect 45502 406658 45586 406894
rect 45822 406658 45854 406894
rect 45234 406574 45854 406658
rect 45234 406338 45266 406574
rect 45502 406338 45586 406574
rect 45822 406338 45854 406574
rect 45234 370894 45854 406338
rect 45234 370658 45266 370894
rect 45502 370658 45586 370894
rect 45822 370658 45854 370894
rect 45234 370574 45854 370658
rect 45234 370338 45266 370574
rect 45502 370338 45586 370574
rect 45822 370338 45854 370574
rect 45234 334894 45854 370338
rect 45234 334658 45266 334894
rect 45502 334658 45586 334894
rect 45822 334658 45854 334894
rect 45234 334574 45854 334658
rect 45234 334338 45266 334574
rect 45502 334338 45586 334574
rect 45822 334338 45854 334574
rect 45234 298894 45854 334338
rect 45234 298658 45266 298894
rect 45502 298658 45586 298894
rect 45822 298658 45854 298894
rect 45234 298574 45854 298658
rect 45234 298338 45266 298574
rect 45502 298338 45586 298574
rect 45822 298338 45854 298574
rect 45234 262894 45854 298338
rect 45234 262658 45266 262894
rect 45502 262658 45586 262894
rect 45822 262658 45854 262894
rect 45234 262574 45854 262658
rect 45234 262338 45266 262574
rect 45502 262338 45586 262574
rect 45822 262338 45854 262574
rect 45234 226894 45854 262338
rect 45234 226658 45266 226894
rect 45502 226658 45586 226894
rect 45822 226658 45854 226894
rect 45234 226574 45854 226658
rect 45234 226338 45266 226574
rect 45502 226338 45586 226574
rect 45822 226338 45854 226574
rect 45234 190894 45854 226338
rect 45234 190658 45266 190894
rect 45502 190658 45586 190894
rect 45822 190658 45854 190894
rect 45234 190574 45854 190658
rect 45234 190338 45266 190574
rect 45502 190338 45586 190574
rect 45822 190338 45854 190574
rect 45234 154894 45854 190338
rect 45234 154658 45266 154894
rect 45502 154658 45586 154894
rect 45822 154658 45854 154894
rect 45234 154574 45854 154658
rect 45234 154338 45266 154574
rect 45502 154338 45586 154574
rect 45822 154338 45854 154574
rect 45234 118894 45854 154338
rect 45234 118658 45266 118894
rect 45502 118658 45586 118894
rect 45822 118658 45854 118894
rect 45234 118574 45854 118658
rect 45234 118338 45266 118574
rect 45502 118338 45586 118574
rect 45822 118338 45854 118574
rect 45234 82894 45854 118338
rect 45234 82658 45266 82894
rect 45502 82658 45586 82894
rect 45822 82658 45854 82894
rect 45234 82574 45854 82658
rect 45234 82338 45266 82574
rect 45502 82338 45586 82574
rect 45822 82338 45854 82574
rect 45234 46894 45854 82338
rect 45234 46658 45266 46894
rect 45502 46658 45586 46894
rect 45822 46658 45854 46894
rect 45234 46574 45854 46658
rect 45234 46338 45266 46574
rect 45502 46338 45586 46574
rect 45822 46338 45854 46574
rect 45234 10894 45854 46338
rect 45234 10658 45266 10894
rect 45502 10658 45586 10894
rect 45822 10658 45854 10894
rect 45234 10574 45854 10658
rect 45234 10338 45266 10574
rect 45502 10338 45586 10574
rect 45822 10338 45854 10574
rect 45234 -4186 45854 10338
rect 45234 -4422 45266 -4186
rect 45502 -4422 45586 -4186
rect 45822 -4422 45854 -4186
rect 45234 -4506 45854 -4422
rect 45234 -4742 45266 -4506
rect 45502 -4742 45586 -4506
rect 45822 -4742 45854 -4506
rect 45234 -5734 45854 -4742
rect 48954 698614 49574 710042
rect 66954 711558 67574 711590
rect 66954 711322 66986 711558
rect 67222 711322 67306 711558
rect 67542 711322 67574 711558
rect 66954 711238 67574 711322
rect 66954 711002 66986 711238
rect 67222 711002 67306 711238
rect 67542 711002 67574 711238
rect 63234 709638 63854 709670
rect 63234 709402 63266 709638
rect 63502 709402 63586 709638
rect 63822 709402 63854 709638
rect 63234 709318 63854 709402
rect 63234 709082 63266 709318
rect 63502 709082 63586 709318
rect 63822 709082 63854 709318
rect 59514 707718 60134 707750
rect 59514 707482 59546 707718
rect 59782 707482 59866 707718
rect 60102 707482 60134 707718
rect 59514 707398 60134 707482
rect 59514 707162 59546 707398
rect 59782 707162 59866 707398
rect 60102 707162 60134 707398
rect 48954 698378 48986 698614
rect 49222 698378 49306 698614
rect 49542 698378 49574 698614
rect 48954 698294 49574 698378
rect 48954 698058 48986 698294
rect 49222 698058 49306 698294
rect 49542 698058 49574 698294
rect 48954 662614 49574 698058
rect 48954 662378 48986 662614
rect 49222 662378 49306 662614
rect 49542 662378 49574 662614
rect 48954 662294 49574 662378
rect 48954 662058 48986 662294
rect 49222 662058 49306 662294
rect 49542 662058 49574 662294
rect 48954 626614 49574 662058
rect 48954 626378 48986 626614
rect 49222 626378 49306 626614
rect 49542 626378 49574 626614
rect 48954 626294 49574 626378
rect 48954 626058 48986 626294
rect 49222 626058 49306 626294
rect 49542 626058 49574 626294
rect 48954 590614 49574 626058
rect 48954 590378 48986 590614
rect 49222 590378 49306 590614
rect 49542 590378 49574 590614
rect 48954 590294 49574 590378
rect 48954 590058 48986 590294
rect 49222 590058 49306 590294
rect 49542 590058 49574 590294
rect 48954 554614 49574 590058
rect 48954 554378 48986 554614
rect 49222 554378 49306 554614
rect 49542 554378 49574 554614
rect 48954 554294 49574 554378
rect 48954 554058 48986 554294
rect 49222 554058 49306 554294
rect 49542 554058 49574 554294
rect 48954 518614 49574 554058
rect 48954 518378 48986 518614
rect 49222 518378 49306 518614
rect 49542 518378 49574 518614
rect 48954 518294 49574 518378
rect 48954 518058 48986 518294
rect 49222 518058 49306 518294
rect 49542 518058 49574 518294
rect 48954 482614 49574 518058
rect 48954 482378 48986 482614
rect 49222 482378 49306 482614
rect 49542 482378 49574 482614
rect 48954 482294 49574 482378
rect 48954 482058 48986 482294
rect 49222 482058 49306 482294
rect 49542 482058 49574 482294
rect 48954 446614 49574 482058
rect 48954 446378 48986 446614
rect 49222 446378 49306 446614
rect 49542 446378 49574 446614
rect 48954 446294 49574 446378
rect 48954 446058 48986 446294
rect 49222 446058 49306 446294
rect 49542 446058 49574 446294
rect 48954 410614 49574 446058
rect 48954 410378 48986 410614
rect 49222 410378 49306 410614
rect 49542 410378 49574 410614
rect 48954 410294 49574 410378
rect 48954 410058 48986 410294
rect 49222 410058 49306 410294
rect 49542 410058 49574 410294
rect 48954 374614 49574 410058
rect 48954 374378 48986 374614
rect 49222 374378 49306 374614
rect 49542 374378 49574 374614
rect 48954 374294 49574 374378
rect 48954 374058 48986 374294
rect 49222 374058 49306 374294
rect 49542 374058 49574 374294
rect 48954 338614 49574 374058
rect 48954 338378 48986 338614
rect 49222 338378 49306 338614
rect 49542 338378 49574 338614
rect 48954 338294 49574 338378
rect 48954 338058 48986 338294
rect 49222 338058 49306 338294
rect 49542 338058 49574 338294
rect 48954 302614 49574 338058
rect 48954 302378 48986 302614
rect 49222 302378 49306 302614
rect 49542 302378 49574 302614
rect 48954 302294 49574 302378
rect 48954 302058 48986 302294
rect 49222 302058 49306 302294
rect 49542 302058 49574 302294
rect 48954 266614 49574 302058
rect 48954 266378 48986 266614
rect 49222 266378 49306 266614
rect 49542 266378 49574 266614
rect 48954 266294 49574 266378
rect 48954 266058 48986 266294
rect 49222 266058 49306 266294
rect 49542 266058 49574 266294
rect 48954 230614 49574 266058
rect 48954 230378 48986 230614
rect 49222 230378 49306 230614
rect 49542 230378 49574 230614
rect 48954 230294 49574 230378
rect 48954 230058 48986 230294
rect 49222 230058 49306 230294
rect 49542 230058 49574 230294
rect 48954 194614 49574 230058
rect 48954 194378 48986 194614
rect 49222 194378 49306 194614
rect 49542 194378 49574 194614
rect 48954 194294 49574 194378
rect 48954 194058 48986 194294
rect 49222 194058 49306 194294
rect 49542 194058 49574 194294
rect 48954 158614 49574 194058
rect 48954 158378 48986 158614
rect 49222 158378 49306 158614
rect 49542 158378 49574 158614
rect 48954 158294 49574 158378
rect 48954 158058 48986 158294
rect 49222 158058 49306 158294
rect 49542 158058 49574 158294
rect 48954 122614 49574 158058
rect 48954 122378 48986 122614
rect 49222 122378 49306 122614
rect 49542 122378 49574 122614
rect 48954 122294 49574 122378
rect 48954 122058 48986 122294
rect 49222 122058 49306 122294
rect 49542 122058 49574 122294
rect 48954 86614 49574 122058
rect 48954 86378 48986 86614
rect 49222 86378 49306 86614
rect 49542 86378 49574 86614
rect 48954 86294 49574 86378
rect 48954 86058 48986 86294
rect 49222 86058 49306 86294
rect 49542 86058 49574 86294
rect 48954 50614 49574 86058
rect 48954 50378 48986 50614
rect 49222 50378 49306 50614
rect 49542 50378 49574 50614
rect 48954 50294 49574 50378
rect 48954 50058 48986 50294
rect 49222 50058 49306 50294
rect 49542 50058 49574 50294
rect 48954 14614 49574 50058
rect 48954 14378 48986 14614
rect 49222 14378 49306 14614
rect 49542 14378 49574 14614
rect 48954 14294 49574 14378
rect 48954 14058 48986 14294
rect 49222 14058 49306 14294
rect 49542 14058 49574 14294
rect 30954 -7302 30986 -7066
rect 31222 -7302 31306 -7066
rect 31542 -7302 31574 -7066
rect 30954 -7386 31574 -7302
rect 30954 -7622 30986 -7386
rect 31222 -7622 31306 -7386
rect 31542 -7622 31574 -7386
rect 30954 -7654 31574 -7622
rect 48954 -6106 49574 14058
rect 55794 705798 56414 705830
rect 55794 705562 55826 705798
rect 56062 705562 56146 705798
rect 56382 705562 56414 705798
rect 55794 705478 56414 705562
rect 55794 705242 55826 705478
rect 56062 705242 56146 705478
rect 56382 705242 56414 705478
rect 55794 669454 56414 705242
rect 55794 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 56414 669454
rect 55794 669134 56414 669218
rect 55794 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 56414 669134
rect 55794 633454 56414 668898
rect 55794 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 56414 633454
rect 55794 633134 56414 633218
rect 55794 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 56414 633134
rect 55794 597454 56414 632898
rect 55794 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 56414 597454
rect 55794 597134 56414 597218
rect 55794 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 56414 597134
rect 55794 561454 56414 596898
rect 55794 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 56414 561454
rect 55794 561134 56414 561218
rect 55794 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 56414 561134
rect 55794 525454 56414 560898
rect 55794 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 56414 525454
rect 55794 525134 56414 525218
rect 55794 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 56414 525134
rect 55794 489454 56414 524898
rect 55794 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 56414 489454
rect 55794 489134 56414 489218
rect 55794 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 56414 489134
rect 55794 453454 56414 488898
rect 55794 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 56414 453454
rect 55794 453134 56414 453218
rect 55794 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 56414 453134
rect 55794 417454 56414 452898
rect 55794 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 56414 417454
rect 55794 417134 56414 417218
rect 55794 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 56414 417134
rect 55794 381454 56414 416898
rect 55794 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 56414 381454
rect 55794 381134 56414 381218
rect 55794 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 56414 381134
rect 55794 345454 56414 380898
rect 55794 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 56414 345454
rect 55794 345134 56414 345218
rect 55794 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 56414 345134
rect 55794 309454 56414 344898
rect 55794 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 56414 309454
rect 55794 309134 56414 309218
rect 55794 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 56414 309134
rect 55794 273454 56414 308898
rect 55794 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 56414 273454
rect 55794 273134 56414 273218
rect 55794 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 56414 273134
rect 55794 237454 56414 272898
rect 55794 237218 55826 237454
rect 56062 237218 56146 237454
rect 56382 237218 56414 237454
rect 55794 237134 56414 237218
rect 55794 236898 55826 237134
rect 56062 236898 56146 237134
rect 56382 236898 56414 237134
rect 55794 201454 56414 236898
rect 55794 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 56414 201454
rect 55794 201134 56414 201218
rect 55794 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 56414 201134
rect 55794 165454 56414 200898
rect 55794 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 56414 165454
rect 55794 165134 56414 165218
rect 55794 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 56414 165134
rect 55794 129454 56414 164898
rect 55794 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 56414 129454
rect 55794 129134 56414 129218
rect 55794 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 56414 129134
rect 55794 93454 56414 128898
rect 55794 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 56414 93454
rect 55794 93134 56414 93218
rect 55794 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 56414 93134
rect 55794 57454 56414 92898
rect 55794 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 56414 57454
rect 55794 57134 56414 57218
rect 55794 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 56414 57134
rect 55794 21454 56414 56898
rect 55794 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 56414 21454
rect 55794 21134 56414 21218
rect 55794 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 56414 21134
rect 55794 -1306 56414 20898
rect 55794 -1542 55826 -1306
rect 56062 -1542 56146 -1306
rect 56382 -1542 56414 -1306
rect 55794 -1626 56414 -1542
rect 55794 -1862 55826 -1626
rect 56062 -1862 56146 -1626
rect 56382 -1862 56414 -1626
rect 55794 -1894 56414 -1862
rect 59514 673174 60134 707162
rect 59514 672938 59546 673174
rect 59782 672938 59866 673174
rect 60102 672938 60134 673174
rect 59514 672854 60134 672938
rect 59514 672618 59546 672854
rect 59782 672618 59866 672854
rect 60102 672618 60134 672854
rect 59514 637174 60134 672618
rect 59514 636938 59546 637174
rect 59782 636938 59866 637174
rect 60102 636938 60134 637174
rect 59514 636854 60134 636938
rect 59514 636618 59546 636854
rect 59782 636618 59866 636854
rect 60102 636618 60134 636854
rect 59514 601174 60134 636618
rect 59514 600938 59546 601174
rect 59782 600938 59866 601174
rect 60102 600938 60134 601174
rect 59514 600854 60134 600938
rect 59514 600618 59546 600854
rect 59782 600618 59866 600854
rect 60102 600618 60134 600854
rect 59514 565174 60134 600618
rect 59514 564938 59546 565174
rect 59782 564938 59866 565174
rect 60102 564938 60134 565174
rect 59514 564854 60134 564938
rect 59514 564618 59546 564854
rect 59782 564618 59866 564854
rect 60102 564618 60134 564854
rect 59514 529174 60134 564618
rect 59514 528938 59546 529174
rect 59782 528938 59866 529174
rect 60102 528938 60134 529174
rect 59514 528854 60134 528938
rect 59514 528618 59546 528854
rect 59782 528618 59866 528854
rect 60102 528618 60134 528854
rect 59514 493174 60134 528618
rect 59514 492938 59546 493174
rect 59782 492938 59866 493174
rect 60102 492938 60134 493174
rect 59514 492854 60134 492938
rect 59514 492618 59546 492854
rect 59782 492618 59866 492854
rect 60102 492618 60134 492854
rect 59514 457174 60134 492618
rect 59514 456938 59546 457174
rect 59782 456938 59866 457174
rect 60102 456938 60134 457174
rect 59514 456854 60134 456938
rect 59514 456618 59546 456854
rect 59782 456618 59866 456854
rect 60102 456618 60134 456854
rect 59514 421174 60134 456618
rect 59514 420938 59546 421174
rect 59782 420938 59866 421174
rect 60102 420938 60134 421174
rect 59514 420854 60134 420938
rect 59514 420618 59546 420854
rect 59782 420618 59866 420854
rect 60102 420618 60134 420854
rect 59514 385174 60134 420618
rect 59514 384938 59546 385174
rect 59782 384938 59866 385174
rect 60102 384938 60134 385174
rect 59514 384854 60134 384938
rect 59514 384618 59546 384854
rect 59782 384618 59866 384854
rect 60102 384618 60134 384854
rect 59514 349174 60134 384618
rect 59514 348938 59546 349174
rect 59782 348938 59866 349174
rect 60102 348938 60134 349174
rect 59514 348854 60134 348938
rect 59514 348618 59546 348854
rect 59782 348618 59866 348854
rect 60102 348618 60134 348854
rect 59514 313174 60134 348618
rect 59514 312938 59546 313174
rect 59782 312938 59866 313174
rect 60102 312938 60134 313174
rect 59514 312854 60134 312938
rect 59514 312618 59546 312854
rect 59782 312618 59866 312854
rect 60102 312618 60134 312854
rect 59514 277174 60134 312618
rect 59514 276938 59546 277174
rect 59782 276938 59866 277174
rect 60102 276938 60134 277174
rect 59514 276854 60134 276938
rect 59514 276618 59546 276854
rect 59782 276618 59866 276854
rect 60102 276618 60134 276854
rect 59514 241174 60134 276618
rect 59514 240938 59546 241174
rect 59782 240938 59866 241174
rect 60102 240938 60134 241174
rect 59514 240854 60134 240938
rect 59514 240618 59546 240854
rect 59782 240618 59866 240854
rect 60102 240618 60134 240854
rect 59514 205174 60134 240618
rect 59514 204938 59546 205174
rect 59782 204938 59866 205174
rect 60102 204938 60134 205174
rect 59514 204854 60134 204938
rect 59514 204618 59546 204854
rect 59782 204618 59866 204854
rect 60102 204618 60134 204854
rect 59514 169174 60134 204618
rect 59514 168938 59546 169174
rect 59782 168938 59866 169174
rect 60102 168938 60134 169174
rect 59514 168854 60134 168938
rect 59514 168618 59546 168854
rect 59782 168618 59866 168854
rect 60102 168618 60134 168854
rect 59514 133174 60134 168618
rect 59514 132938 59546 133174
rect 59782 132938 59866 133174
rect 60102 132938 60134 133174
rect 59514 132854 60134 132938
rect 59514 132618 59546 132854
rect 59782 132618 59866 132854
rect 60102 132618 60134 132854
rect 59514 97174 60134 132618
rect 59514 96938 59546 97174
rect 59782 96938 59866 97174
rect 60102 96938 60134 97174
rect 59514 96854 60134 96938
rect 59514 96618 59546 96854
rect 59782 96618 59866 96854
rect 60102 96618 60134 96854
rect 59514 61174 60134 96618
rect 59514 60938 59546 61174
rect 59782 60938 59866 61174
rect 60102 60938 60134 61174
rect 59514 60854 60134 60938
rect 59514 60618 59546 60854
rect 59782 60618 59866 60854
rect 60102 60618 60134 60854
rect 59514 25174 60134 60618
rect 59514 24938 59546 25174
rect 59782 24938 59866 25174
rect 60102 24938 60134 25174
rect 59514 24854 60134 24938
rect 59514 24618 59546 24854
rect 59782 24618 59866 24854
rect 60102 24618 60134 24854
rect 59514 -3226 60134 24618
rect 59514 -3462 59546 -3226
rect 59782 -3462 59866 -3226
rect 60102 -3462 60134 -3226
rect 59514 -3546 60134 -3462
rect 59514 -3782 59546 -3546
rect 59782 -3782 59866 -3546
rect 60102 -3782 60134 -3546
rect 59514 -3814 60134 -3782
rect 63234 676894 63854 709082
rect 63234 676658 63266 676894
rect 63502 676658 63586 676894
rect 63822 676658 63854 676894
rect 63234 676574 63854 676658
rect 63234 676338 63266 676574
rect 63502 676338 63586 676574
rect 63822 676338 63854 676574
rect 63234 640894 63854 676338
rect 63234 640658 63266 640894
rect 63502 640658 63586 640894
rect 63822 640658 63854 640894
rect 63234 640574 63854 640658
rect 63234 640338 63266 640574
rect 63502 640338 63586 640574
rect 63822 640338 63854 640574
rect 63234 604894 63854 640338
rect 63234 604658 63266 604894
rect 63502 604658 63586 604894
rect 63822 604658 63854 604894
rect 63234 604574 63854 604658
rect 63234 604338 63266 604574
rect 63502 604338 63586 604574
rect 63822 604338 63854 604574
rect 63234 568894 63854 604338
rect 63234 568658 63266 568894
rect 63502 568658 63586 568894
rect 63822 568658 63854 568894
rect 63234 568574 63854 568658
rect 63234 568338 63266 568574
rect 63502 568338 63586 568574
rect 63822 568338 63854 568574
rect 63234 532894 63854 568338
rect 63234 532658 63266 532894
rect 63502 532658 63586 532894
rect 63822 532658 63854 532894
rect 63234 532574 63854 532658
rect 63234 532338 63266 532574
rect 63502 532338 63586 532574
rect 63822 532338 63854 532574
rect 63234 496894 63854 532338
rect 63234 496658 63266 496894
rect 63502 496658 63586 496894
rect 63822 496658 63854 496894
rect 63234 496574 63854 496658
rect 63234 496338 63266 496574
rect 63502 496338 63586 496574
rect 63822 496338 63854 496574
rect 63234 460894 63854 496338
rect 63234 460658 63266 460894
rect 63502 460658 63586 460894
rect 63822 460658 63854 460894
rect 63234 460574 63854 460658
rect 63234 460338 63266 460574
rect 63502 460338 63586 460574
rect 63822 460338 63854 460574
rect 63234 424894 63854 460338
rect 63234 424658 63266 424894
rect 63502 424658 63586 424894
rect 63822 424658 63854 424894
rect 63234 424574 63854 424658
rect 63234 424338 63266 424574
rect 63502 424338 63586 424574
rect 63822 424338 63854 424574
rect 63234 388894 63854 424338
rect 63234 388658 63266 388894
rect 63502 388658 63586 388894
rect 63822 388658 63854 388894
rect 63234 388574 63854 388658
rect 63234 388338 63266 388574
rect 63502 388338 63586 388574
rect 63822 388338 63854 388574
rect 63234 352894 63854 388338
rect 63234 352658 63266 352894
rect 63502 352658 63586 352894
rect 63822 352658 63854 352894
rect 63234 352574 63854 352658
rect 63234 352338 63266 352574
rect 63502 352338 63586 352574
rect 63822 352338 63854 352574
rect 63234 316894 63854 352338
rect 63234 316658 63266 316894
rect 63502 316658 63586 316894
rect 63822 316658 63854 316894
rect 63234 316574 63854 316658
rect 63234 316338 63266 316574
rect 63502 316338 63586 316574
rect 63822 316338 63854 316574
rect 63234 280894 63854 316338
rect 63234 280658 63266 280894
rect 63502 280658 63586 280894
rect 63822 280658 63854 280894
rect 63234 280574 63854 280658
rect 63234 280338 63266 280574
rect 63502 280338 63586 280574
rect 63822 280338 63854 280574
rect 63234 244894 63854 280338
rect 63234 244658 63266 244894
rect 63502 244658 63586 244894
rect 63822 244658 63854 244894
rect 63234 244574 63854 244658
rect 63234 244338 63266 244574
rect 63502 244338 63586 244574
rect 63822 244338 63854 244574
rect 63234 208894 63854 244338
rect 63234 208658 63266 208894
rect 63502 208658 63586 208894
rect 63822 208658 63854 208894
rect 63234 208574 63854 208658
rect 63234 208338 63266 208574
rect 63502 208338 63586 208574
rect 63822 208338 63854 208574
rect 63234 172894 63854 208338
rect 63234 172658 63266 172894
rect 63502 172658 63586 172894
rect 63822 172658 63854 172894
rect 63234 172574 63854 172658
rect 63234 172338 63266 172574
rect 63502 172338 63586 172574
rect 63822 172338 63854 172574
rect 63234 136894 63854 172338
rect 63234 136658 63266 136894
rect 63502 136658 63586 136894
rect 63822 136658 63854 136894
rect 63234 136574 63854 136658
rect 63234 136338 63266 136574
rect 63502 136338 63586 136574
rect 63822 136338 63854 136574
rect 63234 100894 63854 136338
rect 63234 100658 63266 100894
rect 63502 100658 63586 100894
rect 63822 100658 63854 100894
rect 63234 100574 63854 100658
rect 63234 100338 63266 100574
rect 63502 100338 63586 100574
rect 63822 100338 63854 100574
rect 63234 64894 63854 100338
rect 63234 64658 63266 64894
rect 63502 64658 63586 64894
rect 63822 64658 63854 64894
rect 63234 64574 63854 64658
rect 63234 64338 63266 64574
rect 63502 64338 63586 64574
rect 63822 64338 63854 64574
rect 63234 28894 63854 64338
rect 63234 28658 63266 28894
rect 63502 28658 63586 28894
rect 63822 28658 63854 28894
rect 63234 28574 63854 28658
rect 63234 28338 63266 28574
rect 63502 28338 63586 28574
rect 63822 28338 63854 28574
rect 63234 -5146 63854 28338
rect 63234 -5382 63266 -5146
rect 63502 -5382 63586 -5146
rect 63822 -5382 63854 -5146
rect 63234 -5466 63854 -5382
rect 63234 -5702 63266 -5466
rect 63502 -5702 63586 -5466
rect 63822 -5702 63854 -5466
rect 63234 -5734 63854 -5702
rect 66954 680614 67574 711002
rect 84954 710598 85574 711590
rect 84954 710362 84986 710598
rect 85222 710362 85306 710598
rect 85542 710362 85574 710598
rect 84954 710278 85574 710362
rect 84954 710042 84986 710278
rect 85222 710042 85306 710278
rect 85542 710042 85574 710278
rect 81234 708678 81854 709670
rect 81234 708442 81266 708678
rect 81502 708442 81586 708678
rect 81822 708442 81854 708678
rect 81234 708358 81854 708442
rect 81234 708122 81266 708358
rect 81502 708122 81586 708358
rect 81822 708122 81854 708358
rect 77514 706758 78134 707750
rect 77514 706522 77546 706758
rect 77782 706522 77866 706758
rect 78102 706522 78134 706758
rect 77514 706438 78134 706522
rect 77514 706202 77546 706438
rect 77782 706202 77866 706438
rect 78102 706202 78134 706438
rect 66954 680378 66986 680614
rect 67222 680378 67306 680614
rect 67542 680378 67574 680614
rect 66954 680294 67574 680378
rect 66954 680058 66986 680294
rect 67222 680058 67306 680294
rect 67542 680058 67574 680294
rect 66954 644614 67574 680058
rect 66954 644378 66986 644614
rect 67222 644378 67306 644614
rect 67542 644378 67574 644614
rect 66954 644294 67574 644378
rect 66954 644058 66986 644294
rect 67222 644058 67306 644294
rect 67542 644058 67574 644294
rect 66954 608614 67574 644058
rect 66954 608378 66986 608614
rect 67222 608378 67306 608614
rect 67542 608378 67574 608614
rect 66954 608294 67574 608378
rect 66954 608058 66986 608294
rect 67222 608058 67306 608294
rect 67542 608058 67574 608294
rect 66954 572614 67574 608058
rect 66954 572378 66986 572614
rect 67222 572378 67306 572614
rect 67542 572378 67574 572614
rect 66954 572294 67574 572378
rect 66954 572058 66986 572294
rect 67222 572058 67306 572294
rect 67542 572058 67574 572294
rect 66954 536614 67574 572058
rect 66954 536378 66986 536614
rect 67222 536378 67306 536614
rect 67542 536378 67574 536614
rect 66954 536294 67574 536378
rect 66954 536058 66986 536294
rect 67222 536058 67306 536294
rect 67542 536058 67574 536294
rect 66954 500614 67574 536058
rect 66954 500378 66986 500614
rect 67222 500378 67306 500614
rect 67542 500378 67574 500614
rect 66954 500294 67574 500378
rect 66954 500058 66986 500294
rect 67222 500058 67306 500294
rect 67542 500058 67574 500294
rect 66954 464614 67574 500058
rect 66954 464378 66986 464614
rect 67222 464378 67306 464614
rect 67542 464378 67574 464614
rect 66954 464294 67574 464378
rect 66954 464058 66986 464294
rect 67222 464058 67306 464294
rect 67542 464058 67574 464294
rect 66954 428614 67574 464058
rect 66954 428378 66986 428614
rect 67222 428378 67306 428614
rect 67542 428378 67574 428614
rect 66954 428294 67574 428378
rect 66954 428058 66986 428294
rect 67222 428058 67306 428294
rect 67542 428058 67574 428294
rect 66954 392614 67574 428058
rect 66954 392378 66986 392614
rect 67222 392378 67306 392614
rect 67542 392378 67574 392614
rect 66954 392294 67574 392378
rect 66954 392058 66986 392294
rect 67222 392058 67306 392294
rect 67542 392058 67574 392294
rect 66954 356614 67574 392058
rect 66954 356378 66986 356614
rect 67222 356378 67306 356614
rect 67542 356378 67574 356614
rect 66954 356294 67574 356378
rect 66954 356058 66986 356294
rect 67222 356058 67306 356294
rect 67542 356058 67574 356294
rect 66954 320614 67574 356058
rect 66954 320378 66986 320614
rect 67222 320378 67306 320614
rect 67542 320378 67574 320614
rect 66954 320294 67574 320378
rect 66954 320058 66986 320294
rect 67222 320058 67306 320294
rect 67542 320058 67574 320294
rect 66954 284614 67574 320058
rect 66954 284378 66986 284614
rect 67222 284378 67306 284614
rect 67542 284378 67574 284614
rect 66954 284294 67574 284378
rect 66954 284058 66986 284294
rect 67222 284058 67306 284294
rect 67542 284058 67574 284294
rect 66954 248614 67574 284058
rect 66954 248378 66986 248614
rect 67222 248378 67306 248614
rect 67542 248378 67574 248614
rect 66954 248294 67574 248378
rect 66954 248058 66986 248294
rect 67222 248058 67306 248294
rect 67542 248058 67574 248294
rect 66954 212614 67574 248058
rect 66954 212378 66986 212614
rect 67222 212378 67306 212614
rect 67542 212378 67574 212614
rect 66954 212294 67574 212378
rect 66954 212058 66986 212294
rect 67222 212058 67306 212294
rect 67542 212058 67574 212294
rect 66954 176614 67574 212058
rect 66954 176378 66986 176614
rect 67222 176378 67306 176614
rect 67542 176378 67574 176614
rect 66954 176294 67574 176378
rect 66954 176058 66986 176294
rect 67222 176058 67306 176294
rect 67542 176058 67574 176294
rect 66954 140614 67574 176058
rect 66954 140378 66986 140614
rect 67222 140378 67306 140614
rect 67542 140378 67574 140614
rect 66954 140294 67574 140378
rect 66954 140058 66986 140294
rect 67222 140058 67306 140294
rect 67542 140058 67574 140294
rect 66954 104614 67574 140058
rect 66954 104378 66986 104614
rect 67222 104378 67306 104614
rect 67542 104378 67574 104614
rect 66954 104294 67574 104378
rect 66954 104058 66986 104294
rect 67222 104058 67306 104294
rect 67542 104058 67574 104294
rect 66954 68614 67574 104058
rect 66954 68378 66986 68614
rect 67222 68378 67306 68614
rect 67542 68378 67574 68614
rect 66954 68294 67574 68378
rect 66954 68058 66986 68294
rect 67222 68058 67306 68294
rect 67542 68058 67574 68294
rect 66954 32614 67574 68058
rect 66954 32378 66986 32614
rect 67222 32378 67306 32614
rect 67542 32378 67574 32614
rect 66954 32294 67574 32378
rect 66954 32058 66986 32294
rect 67222 32058 67306 32294
rect 67542 32058 67574 32294
rect 48954 -6342 48986 -6106
rect 49222 -6342 49306 -6106
rect 49542 -6342 49574 -6106
rect 48954 -6426 49574 -6342
rect 48954 -6662 48986 -6426
rect 49222 -6662 49306 -6426
rect 49542 -6662 49574 -6426
rect 48954 -7654 49574 -6662
rect 66954 -7066 67574 32058
rect 73794 704838 74414 705830
rect 73794 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 74414 704838
rect 73794 704518 74414 704602
rect 73794 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 74414 704518
rect 73794 687454 74414 704282
rect 73794 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 74414 687454
rect 73794 687134 74414 687218
rect 73794 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 74414 687134
rect 73794 651454 74414 686898
rect 73794 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 74414 651454
rect 73794 651134 74414 651218
rect 73794 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 74414 651134
rect 73794 615454 74414 650898
rect 73794 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 74414 615454
rect 73794 615134 74414 615218
rect 73794 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 74414 615134
rect 73794 579454 74414 614898
rect 73794 579218 73826 579454
rect 74062 579218 74146 579454
rect 74382 579218 74414 579454
rect 73794 579134 74414 579218
rect 73794 578898 73826 579134
rect 74062 578898 74146 579134
rect 74382 578898 74414 579134
rect 73794 543454 74414 578898
rect 73794 543218 73826 543454
rect 74062 543218 74146 543454
rect 74382 543218 74414 543454
rect 73794 543134 74414 543218
rect 73794 542898 73826 543134
rect 74062 542898 74146 543134
rect 74382 542898 74414 543134
rect 73794 507454 74414 542898
rect 73794 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 74414 507454
rect 73794 507134 74414 507218
rect 73794 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 74414 507134
rect 73794 471454 74414 506898
rect 73794 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 74414 471454
rect 73794 471134 74414 471218
rect 73794 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 74414 471134
rect 73794 435454 74414 470898
rect 73794 435218 73826 435454
rect 74062 435218 74146 435454
rect 74382 435218 74414 435454
rect 73794 435134 74414 435218
rect 73794 434898 73826 435134
rect 74062 434898 74146 435134
rect 74382 434898 74414 435134
rect 73794 399454 74414 434898
rect 73794 399218 73826 399454
rect 74062 399218 74146 399454
rect 74382 399218 74414 399454
rect 73794 399134 74414 399218
rect 73794 398898 73826 399134
rect 74062 398898 74146 399134
rect 74382 398898 74414 399134
rect 73794 363454 74414 398898
rect 73794 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 74414 363454
rect 73794 363134 74414 363218
rect 73794 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 74414 363134
rect 73794 327454 74414 362898
rect 73794 327218 73826 327454
rect 74062 327218 74146 327454
rect 74382 327218 74414 327454
rect 73794 327134 74414 327218
rect 73794 326898 73826 327134
rect 74062 326898 74146 327134
rect 74382 326898 74414 327134
rect 73794 291454 74414 326898
rect 73794 291218 73826 291454
rect 74062 291218 74146 291454
rect 74382 291218 74414 291454
rect 73794 291134 74414 291218
rect 73794 290898 73826 291134
rect 74062 290898 74146 291134
rect 74382 290898 74414 291134
rect 73794 255454 74414 290898
rect 73794 255218 73826 255454
rect 74062 255218 74146 255454
rect 74382 255218 74414 255454
rect 73794 255134 74414 255218
rect 73794 254898 73826 255134
rect 74062 254898 74146 255134
rect 74382 254898 74414 255134
rect 73794 219454 74414 254898
rect 73794 219218 73826 219454
rect 74062 219218 74146 219454
rect 74382 219218 74414 219454
rect 73794 219134 74414 219218
rect 73794 218898 73826 219134
rect 74062 218898 74146 219134
rect 74382 218898 74414 219134
rect 73794 183454 74414 218898
rect 73794 183218 73826 183454
rect 74062 183218 74146 183454
rect 74382 183218 74414 183454
rect 73794 183134 74414 183218
rect 73794 182898 73826 183134
rect 74062 182898 74146 183134
rect 74382 182898 74414 183134
rect 73794 147454 74414 182898
rect 73794 147218 73826 147454
rect 74062 147218 74146 147454
rect 74382 147218 74414 147454
rect 73794 147134 74414 147218
rect 73794 146898 73826 147134
rect 74062 146898 74146 147134
rect 74382 146898 74414 147134
rect 73794 111454 74414 146898
rect 73794 111218 73826 111454
rect 74062 111218 74146 111454
rect 74382 111218 74414 111454
rect 73794 111134 74414 111218
rect 73794 110898 73826 111134
rect 74062 110898 74146 111134
rect 74382 110898 74414 111134
rect 73794 75454 74414 110898
rect 73794 75218 73826 75454
rect 74062 75218 74146 75454
rect 74382 75218 74414 75454
rect 73794 75134 74414 75218
rect 73794 74898 73826 75134
rect 74062 74898 74146 75134
rect 74382 74898 74414 75134
rect 73794 39454 74414 74898
rect 73794 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 74414 39454
rect 73794 39134 74414 39218
rect 73794 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 74414 39134
rect 73794 3454 74414 38898
rect 73794 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 74414 3454
rect 73794 3134 74414 3218
rect 73794 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 74414 3134
rect 73794 -346 74414 2898
rect 73794 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 74414 -346
rect 73794 -666 74414 -582
rect 73794 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 74414 -666
rect 73794 -1894 74414 -902
rect 77514 691174 78134 706202
rect 77514 690938 77546 691174
rect 77782 690938 77866 691174
rect 78102 690938 78134 691174
rect 77514 690854 78134 690938
rect 77514 690618 77546 690854
rect 77782 690618 77866 690854
rect 78102 690618 78134 690854
rect 77514 655174 78134 690618
rect 77514 654938 77546 655174
rect 77782 654938 77866 655174
rect 78102 654938 78134 655174
rect 77514 654854 78134 654938
rect 77514 654618 77546 654854
rect 77782 654618 77866 654854
rect 78102 654618 78134 654854
rect 77514 619174 78134 654618
rect 77514 618938 77546 619174
rect 77782 618938 77866 619174
rect 78102 618938 78134 619174
rect 77514 618854 78134 618938
rect 77514 618618 77546 618854
rect 77782 618618 77866 618854
rect 78102 618618 78134 618854
rect 77514 583174 78134 618618
rect 77514 582938 77546 583174
rect 77782 582938 77866 583174
rect 78102 582938 78134 583174
rect 77514 582854 78134 582938
rect 77514 582618 77546 582854
rect 77782 582618 77866 582854
rect 78102 582618 78134 582854
rect 77514 547174 78134 582618
rect 77514 546938 77546 547174
rect 77782 546938 77866 547174
rect 78102 546938 78134 547174
rect 77514 546854 78134 546938
rect 77514 546618 77546 546854
rect 77782 546618 77866 546854
rect 78102 546618 78134 546854
rect 77514 511174 78134 546618
rect 77514 510938 77546 511174
rect 77782 510938 77866 511174
rect 78102 510938 78134 511174
rect 77514 510854 78134 510938
rect 77514 510618 77546 510854
rect 77782 510618 77866 510854
rect 78102 510618 78134 510854
rect 77514 475174 78134 510618
rect 77514 474938 77546 475174
rect 77782 474938 77866 475174
rect 78102 474938 78134 475174
rect 77514 474854 78134 474938
rect 77514 474618 77546 474854
rect 77782 474618 77866 474854
rect 78102 474618 78134 474854
rect 77514 439174 78134 474618
rect 77514 438938 77546 439174
rect 77782 438938 77866 439174
rect 78102 438938 78134 439174
rect 77514 438854 78134 438938
rect 77514 438618 77546 438854
rect 77782 438618 77866 438854
rect 78102 438618 78134 438854
rect 77514 403174 78134 438618
rect 77514 402938 77546 403174
rect 77782 402938 77866 403174
rect 78102 402938 78134 403174
rect 77514 402854 78134 402938
rect 77514 402618 77546 402854
rect 77782 402618 77866 402854
rect 78102 402618 78134 402854
rect 77514 367174 78134 402618
rect 77514 366938 77546 367174
rect 77782 366938 77866 367174
rect 78102 366938 78134 367174
rect 77514 366854 78134 366938
rect 77514 366618 77546 366854
rect 77782 366618 77866 366854
rect 78102 366618 78134 366854
rect 77514 331174 78134 366618
rect 77514 330938 77546 331174
rect 77782 330938 77866 331174
rect 78102 330938 78134 331174
rect 77514 330854 78134 330938
rect 77514 330618 77546 330854
rect 77782 330618 77866 330854
rect 78102 330618 78134 330854
rect 77514 295174 78134 330618
rect 77514 294938 77546 295174
rect 77782 294938 77866 295174
rect 78102 294938 78134 295174
rect 77514 294854 78134 294938
rect 77514 294618 77546 294854
rect 77782 294618 77866 294854
rect 78102 294618 78134 294854
rect 77514 259174 78134 294618
rect 77514 258938 77546 259174
rect 77782 258938 77866 259174
rect 78102 258938 78134 259174
rect 77514 258854 78134 258938
rect 77514 258618 77546 258854
rect 77782 258618 77866 258854
rect 78102 258618 78134 258854
rect 77514 223174 78134 258618
rect 77514 222938 77546 223174
rect 77782 222938 77866 223174
rect 78102 222938 78134 223174
rect 77514 222854 78134 222938
rect 77514 222618 77546 222854
rect 77782 222618 77866 222854
rect 78102 222618 78134 222854
rect 77514 187174 78134 222618
rect 77514 186938 77546 187174
rect 77782 186938 77866 187174
rect 78102 186938 78134 187174
rect 77514 186854 78134 186938
rect 77514 186618 77546 186854
rect 77782 186618 77866 186854
rect 78102 186618 78134 186854
rect 77514 151174 78134 186618
rect 77514 150938 77546 151174
rect 77782 150938 77866 151174
rect 78102 150938 78134 151174
rect 77514 150854 78134 150938
rect 77514 150618 77546 150854
rect 77782 150618 77866 150854
rect 78102 150618 78134 150854
rect 77514 115174 78134 150618
rect 77514 114938 77546 115174
rect 77782 114938 77866 115174
rect 78102 114938 78134 115174
rect 77514 114854 78134 114938
rect 77514 114618 77546 114854
rect 77782 114618 77866 114854
rect 78102 114618 78134 114854
rect 77514 79174 78134 114618
rect 77514 78938 77546 79174
rect 77782 78938 77866 79174
rect 78102 78938 78134 79174
rect 77514 78854 78134 78938
rect 77514 78618 77546 78854
rect 77782 78618 77866 78854
rect 78102 78618 78134 78854
rect 77514 43174 78134 78618
rect 77514 42938 77546 43174
rect 77782 42938 77866 43174
rect 78102 42938 78134 43174
rect 77514 42854 78134 42938
rect 77514 42618 77546 42854
rect 77782 42618 77866 42854
rect 78102 42618 78134 42854
rect 77514 7174 78134 42618
rect 77514 6938 77546 7174
rect 77782 6938 77866 7174
rect 78102 6938 78134 7174
rect 77514 6854 78134 6938
rect 77514 6618 77546 6854
rect 77782 6618 77866 6854
rect 78102 6618 78134 6854
rect 77514 -2266 78134 6618
rect 77514 -2502 77546 -2266
rect 77782 -2502 77866 -2266
rect 78102 -2502 78134 -2266
rect 77514 -2586 78134 -2502
rect 77514 -2822 77546 -2586
rect 77782 -2822 77866 -2586
rect 78102 -2822 78134 -2586
rect 77514 -3814 78134 -2822
rect 81234 694894 81854 708122
rect 81234 694658 81266 694894
rect 81502 694658 81586 694894
rect 81822 694658 81854 694894
rect 81234 694574 81854 694658
rect 81234 694338 81266 694574
rect 81502 694338 81586 694574
rect 81822 694338 81854 694574
rect 81234 658894 81854 694338
rect 81234 658658 81266 658894
rect 81502 658658 81586 658894
rect 81822 658658 81854 658894
rect 81234 658574 81854 658658
rect 81234 658338 81266 658574
rect 81502 658338 81586 658574
rect 81822 658338 81854 658574
rect 81234 622894 81854 658338
rect 81234 622658 81266 622894
rect 81502 622658 81586 622894
rect 81822 622658 81854 622894
rect 81234 622574 81854 622658
rect 81234 622338 81266 622574
rect 81502 622338 81586 622574
rect 81822 622338 81854 622574
rect 81234 586894 81854 622338
rect 81234 586658 81266 586894
rect 81502 586658 81586 586894
rect 81822 586658 81854 586894
rect 81234 586574 81854 586658
rect 81234 586338 81266 586574
rect 81502 586338 81586 586574
rect 81822 586338 81854 586574
rect 81234 550894 81854 586338
rect 81234 550658 81266 550894
rect 81502 550658 81586 550894
rect 81822 550658 81854 550894
rect 81234 550574 81854 550658
rect 81234 550338 81266 550574
rect 81502 550338 81586 550574
rect 81822 550338 81854 550574
rect 81234 514894 81854 550338
rect 81234 514658 81266 514894
rect 81502 514658 81586 514894
rect 81822 514658 81854 514894
rect 81234 514574 81854 514658
rect 81234 514338 81266 514574
rect 81502 514338 81586 514574
rect 81822 514338 81854 514574
rect 81234 478894 81854 514338
rect 81234 478658 81266 478894
rect 81502 478658 81586 478894
rect 81822 478658 81854 478894
rect 81234 478574 81854 478658
rect 81234 478338 81266 478574
rect 81502 478338 81586 478574
rect 81822 478338 81854 478574
rect 81234 442894 81854 478338
rect 81234 442658 81266 442894
rect 81502 442658 81586 442894
rect 81822 442658 81854 442894
rect 81234 442574 81854 442658
rect 81234 442338 81266 442574
rect 81502 442338 81586 442574
rect 81822 442338 81854 442574
rect 81234 406894 81854 442338
rect 81234 406658 81266 406894
rect 81502 406658 81586 406894
rect 81822 406658 81854 406894
rect 81234 406574 81854 406658
rect 81234 406338 81266 406574
rect 81502 406338 81586 406574
rect 81822 406338 81854 406574
rect 81234 370894 81854 406338
rect 81234 370658 81266 370894
rect 81502 370658 81586 370894
rect 81822 370658 81854 370894
rect 81234 370574 81854 370658
rect 81234 370338 81266 370574
rect 81502 370338 81586 370574
rect 81822 370338 81854 370574
rect 81234 334894 81854 370338
rect 81234 334658 81266 334894
rect 81502 334658 81586 334894
rect 81822 334658 81854 334894
rect 81234 334574 81854 334658
rect 81234 334338 81266 334574
rect 81502 334338 81586 334574
rect 81822 334338 81854 334574
rect 81234 298894 81854 334338
rect 81234 298658 81266 298894
rect 81502 298658 81586 298894
rect 81822 298658 81854 298894
rect 81234 298574 81854 298658
rect 81234 298338 81266 298574
rect 81502 298338 81586 298574
rect 81822 298338 81854 298574
rect 81234 262894 81854 298338
rect 81234 262658 81266 262894
rect 81502 262658 81586 262894
rect 81822 262658 81854 262894
rect 81234 262574 81854 262658
rect 81234 262338 81266 262574
rect 81502 262338 81586 262574
rect 81822 262338 81854 262574
rect 81234 226894 81854 262338
rect 81234 226658 81266 226894
rect 81502 226658 81586 226894
rect 81822 226658 81854 226894
rect 81234 226574 81854 226658
rect 81234 226338 81266 226574
rect 81502 226338 81586 226574
rect 81822 226338 81854 226574
rect 81234 190894 81854 226338
rect 81234 190658 81266 190894
rect 81502 190658 81586 190894
rect 81822 190658 81854 190894
rect 81234 190574 81854 190658
rect 81234 190338 81266 190574
rect 81502 190338 81586 190574
rect 81822 190338 81854 190574
rect 81234 154894 81854 190338
rect 81234 154658 81266 154894
rect 81502 154658 81586 154894
rect 81822 154658 81854 154894
rect 81234 154574 81854 154658
rect 81234 154338 81266 154574
rect 81502 154338 81586 154574
rect 81822 154338 81854 154574
rect 81234 118894 81854 154338
rect 81234 118658 81266 118894
rect 81502 118658 81586 118894
rect 81822 118658 81854 118894
rect 81234 118574 81854 118658
rect 81234 118338 81266 118574
rect 81502 118338 81586 118574
rect 81822 118338 81854 118574
rect 81234 82894 81854 118338
rect 81234 82658 81266 82894
rect 81502 82658 81586 82894
rect 81822 82658 81854 82894
rect 81234 82574 81854 82658
rect 81234 82338 81266 82574
rect 81502 82338 81586 82574
rect 81822 82338 81854 82574
rect 81234 46894 81854 82338
rect 81234 46658 81266 46894
rect 81502 46658 81586 46894
rect 81822 46658 81854 46894
rect 81234 46574 81854 46658
rect 81234 46338 81266 46574
rect 81502 46338 81586 46574
rect 81822 46338 81854 46574
rect 81234 10894 81854 46338
rect 81234 10658 81266 10894
rect 81502 10658 81586 10894
rect 81822 10658 81854 10894
rect 81234 10574 81854 10658
rect 81234 10338 81266 10574
rect 81502 10338 81586 10574
rect 81822 10338 81854 10574
rect 81234 -4186 81854 10338
rect 81234 -4422 81266 -4186
rect 81502 -4422 81586 -4186
rect 81822 -4422 81854 -4186
rect 81234 -4506 81854 -4422
rect 81234 -4742 81266 -4506
rect 81502 -4742 81586 -4506
rect 81822 -4742 81854 -4506
rect 81234 -5734 81854 -4742
rect 84954 698614 85574 710042
rect 102954 711558 103574 711590
rect 102954 711322 102986 711558
rect 103222 711322 103306 711558
rect 103542 711322 103574 711558
rect 102954 711238 103574 711322
rect 102954 711002 102986 711238
rect 103222 711002 103306 711238
rect 103542 711002 103574 711238
rect 99234 709638 99854 709670
rect 99234 709402 99266 709638
rect 99502 709402 99586 709638
rect 99822 709402 99854 709638
rect 99234 709318 99854 709402
rect 99234 709082 99266 709318
rect 99502 709082 99586 709318
rect 99822 709082 99854 709318
rect 95514 707718 96134 707750
rect 95514 707482 95546 707718
rect 95782 707482 95866 707718
rect 96102 707482 96134 707718
rect 95514 707398 96134 707482
rect 95514 707162 95546 707398
rect 95782 707162 95866 707398
rect 96102 707162 96134 707398
rect 84954 698378 84986 698614
rect 85222 698378 85306 698614
rect 85542 698378 85574 698614
rect 84954 698294 85574 698378
rect 84954 698058 84986 698294
rect 85222 698058 85306 698294
rect 85542 698058 85574 698294
rect 84954 662614 85574 698058
rect 84954 662378 84986 662614
rect 85222 662378 85306 662614
rect 85542 662378 85574 662614
rect 84954 662294 85574 662378
rect 84954 662058 84986 662294
rect 85222 662058 85306 662294
rect 85542 662058 85574 662294
rect 84954 626614 85574 662058
rect 84954 626378 84986 626614
rect 85222 626378 85306 626614
rect 85542 626378 85574 626614
rect 84954 626294 85574 626378
rect 84954 626058 84986 626294
rect 85222 626058 85306 626294
rect 85542 626058 85574 626294
rect 84954 590614 85574 626058
rect 84954 590378 84986 590614
rect 85222 590378 85306 590614
rect 85542 590378 85574 590614
rect 84954 590294 85574 590378
rect 84954 590058 84986 590294
rect 85222 590058 85306 590294
rect 85542 590058 85574 590294
rect 84954 554614 85574 590058
rect 84954 554378 84986 554614
rect 85222 554378 85306 554614
rect 85542 554378 85574 554614
rect 84954 554294 85574 554378
rect 84954 554058 84986 554294
rect 85222 554058 85306 554294
rect 85542 554058 85574 554294
rect 84954 518614 85574 554058
rect 84954 518378 84986 518614
rect 85222 518378 85306 518614
rect 85542 518378 85574 518614
rect 84954 518294 85574 518378
rect 84954 518058 84986 518294
rect 85222 518058 85306 518294
rect 85542 518058 85574 518294
rect 84954 482614 85574 518058
rect 84954 482378 84986 482614
rect 85222 482378 85306 482614
rect 85542 482378 85574 482614
rect 84954 482294 85574 482378
rect 84954 482058 84986 482294
rect 85222 482058 85306 482294
rect 85542 482058 85574 482294
rect 84954 446614 85574 482058
rect 84954 446378 84986 446614
rect 85222 446378 85306 446614
rect 85542 446378 85574 446614
rect 84954 446294 85574 446378
rect 84954 446058 84986 446294
rect 85222 446058 85306 446294
rect 85542 446058 85574 446294
rect 84954 410614 85574 446058
rect 84954 410378 84986 410614
rect 85222 410378 85306 410614
rect 85542 410378 85574 410614
rect 84954 410294 85574 410378
rect 84954 410058 84986 410294
rect 85222 410058 85306 410294
rect 85542 410058 85574 410294
rect 84954 374614 85574 410058
rect 84954 374378 84986 374614
rect 85222 374378 85306 374614
rect 85542 374378 85574 374614
rect 84954 374294 85574 374378
rect 84954 374058 84986 374294
rect 85222 374058 85306 374294
rect 85542 374058 85574 374294
rect 84954 338614 85574 374058
rect 84954 338378 84986 338614
rect 85222 338378 85306 338614
rect 85542 338378 85574 338614
rect 84954 338294 85574 338378
rect 84954 338058 84986 338294
rect 85222 338058 85306 338294
rect 85542 338058 85574 338294
rect 84954 302614 85574 338058
rect 84954 302378 84986 302614
rect 85222 302378 85306 302614
rect 85542 302378 85574 302614
rect 84954 302294 85574 302378
rect 84954 302058 84986 302294
rect 85222 302058 85306 302294
rect 85542 302058 85574 302294
rect 84954 266614 85574 302058
rect 84954 266378 84986 266614
rect 85222 266378 85306 266614
rect 85542 266378 85574 266614
rect 84954 266294 85574 266378
rect 84954 266058 84986 266294
rect 85222 266058 85306 266294
rect 85542 266058 85574 266294
rect 84954 230614 85574 266058
rect 84954 230378 84986 230614
rect 85222 230378 85306 230614
rect 85542 230378 85574 230614
rect 84954 230294 85574 230378
rect 84954 230058 84986 230294
rect 85222 230058 85306 230294
rect 85542 230058 85574 230294
rect 84954 194614 85574 230058
rect 84954 194378 84986 194614
rect 85222 194378 85306 194614
rect 85542 194378 85574 194614
rect 84954 194294 85574 194378
rect 84954 194058 84986 194294
rect 85222 194058 85306 194294
rect 85542 194058 85574 194294
rect 84954 158614 85574 194058
rect 84954 158378 84986 158614
rect 85222 158378 85306 158614
rect 85542 158378 85574 158614
rect 84954 158294 85574 158378
rect 84954 158058 84986 158294
rect 85222 158058 85306 158294
rect 85542 158058 85574 158294
rect 84954 122614 85574 158058
rect 84954 122378 84986 122614
rect 85222 122378 85306 122614
rect 85542 122378 85574 122614
rect 84954 122294 85574 122378
rect 84954 122058 84986 122294
rect 85222 122058 85306 122294
rect 85542 122058 85574 122294
rect 84954 86614 85574 122058
rect 84954 86378 84986 86614
rect 85222 86378 85306 86614
rect 85542 86378 85574 86614
rect 84954 86294 85574 86378
rect 84954 86058 84986 86294
rect 85222 86058 85306 86294
rect 85542 86058 85574 86294
rect 84954 50614 85574 86058
rect 84954 50378 84986 50614
rect 85222 50378 85306 50614
rect 85542 50378 85574 50614
rect 84954 50294 85574 50378
rect 84954 50058 84986 50294
rect 85222 50058 85306 50294
rect 85542 50058 85574 50294
rect 84954 14614 85574 50058
rect 84954 14378 84986 14614
rect 85222 14378 85306 14614
rect 85542 14378 85574 14614
rect 84954 14294 85574 14378
rect 84954 14058 84986 14294
rect 85222 14058 85306 14294
rect 85542 14058 85574 14294
rect 66954 -7302 66986 -7066
rect 67222 -7302 67306 -7066
rect 67542 -7302 67574 -7066
rect 66954 -7386 67574 -7302
rect 66954 -7622 66986 -7386
rect 67222 -7622 67306 -7386
rect 67542 -7622 67574 -7386
rect 66954 -7654 67574 -7622
rect 84954 -6106 85574 14058
rect 91794 705798 92414 705830
rect 91794 705562 91826 705798
rect 92062 705562 92146 705798
rect 92382 705562 92414 705798
rect 91794 705478 92414 705562
rect 91794 705242 91826 705478
rect 92062 705242 92146 705478
rect 92382 705242 92414 705478
rect 91794 669454 92414 705242
rect 91794 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 92414 669454
rect 91794 669134 92414 669218
rect 91794 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 92414 669134
rect 91794 633454 92414 668898
rect 91794 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 92414 633454
rect 91794 633134 92414 633218
rect 91794 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 92414 633134
rect 91794 597454 92414 632898
rect 91794 597218 91826 597454
rect 92062 597218 92146 597454
rect 92382 597218 92414 597454
rect 91794 597134 92414 597218
rect 91794 596898 91826 597134
rect 92062 596898 92146 597134
rect 92382 596898 92414 597134
rect 91794 561454 92414 596898
rect 91794 561218 91826 561454
rect 92062 561218 92146 561454
rect 92382 561218 92414 561454
rect 91794 561134 92414 561218
rect 91794 560898 91826 561134
rect 92062 560898 92146 561134
rect 92382 560898 92414 561134
rect 91794 525454 92414 560898
rect 91794 525218 91826 525454
rect 92062 525218 92146 525454
rect 92382 525218 92414 525454
rect 91794 525134 92414 525218
rect 91794 524898 91826 525134
rect 92062 524898 92146 525134
rect 92382 524898 92414 525134
rect 91794 489454 92414 524898
rect 91794 489218 91826 489454
rect 92062 489218 92146 489454
rect 92382 489218 92414 489454
rect 91794 489134 92414 489218
rect 91794 488898 91826 489134
rect 92062 488898 92146 489134
rect 92382 488898 92414 489134
rect 91794 453454 92414 488898
rect 91794 453218 91826 453454
rect 92062 453218 92146 453454
rect 92382 453218 92414 453454
rect 91794 453134 92414 453218
rect 91794 452898 91826 453134
rect 92062 452898 92146 453134
rect 92382 452898 92414 453134
rect 91794 417454 92414 452898
rect 91794 417218 91826 417454
rect 92062 417218 92146 417454
rect 92382 417218 92414 417454
rect 91794 417134 92414 417218
rect 91794 416898 91826 417134
rect 92062 416898 92146 417134
rect 92382 416898 92414 417134
rect 91794 381454 92414 416898
rect 91794 381218 91826 381454
rect 92062 381218 92146 381454
rect 92382 381218 92414 381454
rect 91794 381134 92414 381218
rect 91794 380898 91826 381134
rect 92062 380898 92146 381134
rect 92382 380898 92414 381134
rect 91794 345454 92414 380898
rect 91794 345218 91826 345454
rect 92062 345218 92146 345454
rect 92382 345218 92414 345454
rect 91794 345134 92414 345218
rect 91794 344898 91826 345134
rect 92062 344898 92146 345134
rect 92382 344898 92414 345134
rect 91794 309454 92414 344898
rect 91794 309218 91826 309454
rect 92062 309218 92146 309454
rect 92382 309218 92414 309454
rect 91794 309134 92414 309218
rect 91794 308898 91826 309134
rect 92062 308898 92146 309134
rect 92382 308898 92414 309134
rect 91794 273454 92414 308898
rect 91794 273218 91826 273454
rect 92062 273218 92146 273454
rect 92382 273218 92414 273454
rect 91794 273134 92414 273218
rect 91794 272898 91826 273134
rect 92062 272898 92146 273134
rect 92382 272898 92414 273134
rect 91794 237454 92414 272898
rect 91794 237218 91826 237454
rect 92062 237218 92146 237454
rect 92382 237218 92414 237454
rect 91794 237134 92414 237218
rect 91794 236898 91826 237134
rect 92062 236898 92146 237134
rect 92382 236898 92414 237134
rect 91794 201454 92414 236898
rect 91794 201218 91826 201454
rect 92062 201218 92146 201454
rect 92382 201218 92414 201454
rect 91794 201134 92414 201218
rect 91794 200898 91826 201134
rect 92062 200898 92146 201134
rect 92382 200898 92414 201134
rect 91794 165454 92414 200898
rect 91794 165218 91826 165454
rect 92062 165218 92146 165454
rect 92382 165218 92414 165454
rect 91794 165134 92414 165218
rect 91794 164898 91826 165134
rect 92062 164898 92146 165134
rect 92382 164898 92414 165134
rect 91794 129454 92414 164898
rect 91794 129218 91826 129454
rect 92062 129218 92146 129454
rect 92382 129218 92414 129454
rect 91794 129134 92414 129218
rect 91794 128898 91826 129134
rect 92062 128898 92146 129134
rect 92382 128898 92414 129134
rect 91794 93454 92414 128898
rect 91794 93218 91826 93454
rect 92062 93218 92146 93454
rect 92382 93218 92414 93454
rect 91794 93134 92414 93218
rect 91794 92898 91826 93134
rect 92062 92898 92146 93134
rect 92382 92898 92414 93134
rect 91794 57454 92414 92898
rect 91794 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 92414 57454
rect 91794 57134 92414 57218
rect 91794 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 92414 57134
rect 91794 21454 92414 56898
rect 91794 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 92414 21454
rect 91794 21134 92414 21218
rect 91794 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 92414 21134
rect 91794 -1306 92414 20898
rect 91794 -1542 91826 -1306
rect 92062 -1542 92146 -1306
rect 92382 -1542 92414 -1306
rect 91794 -1626 92414 -1542
rect 91794 -1862 91826 -1626
rect 92062 -1862 92146 -1626
rect 92382 -1862 92414 -1626
rect 91794 -1894 92414 -1862
rect 95514 673174 96134 707162
rect 95514 672938 95546 673174
rect 95782 672938 95866 673174
rect 96102 672938 96134 673174
rect 95514 672854 96134 672938
rect 95514 672618 95546 672854
rect 95782 672618 95866 672854
rect 96102 672618 96134 672854
rect 95514 637174 96134 672618
rect 95514 636938 95546 637174
rect 95782 636938 95866 637174
rect 96102 636938 96134 637174
rect 95514 636854 96134 636938
rect 95514 636618 95546 636854
rect 95782 636618 95866 636854
rect 96102 636618 96134 636854
rect 95514 601174 96134 636618
rect 95514 600938 95546 601174
rect 95782 600938 95866 601174
rect 96102 600938 96134 601174
rect 95514 600854 96134 600938
rect 95514 600618 95546 600854
rect 95782 600618 95866 600854
rect 96102 600618 96134 600854
rect 95514 565174 96134 600618
rect 95514 564938 95546 565174
rect 95782 564938 95866 565174
rect 96102 564938 96134 565174
rect 95514 564854 96134 564938
rect 95514 564618 95546 564854
rect 95782 564618 95866 564854
rect 96102 564618 96134 564854
rect 95514 529174 96134 564618
rect 95514 528938 95546 529174
rect 95782 528938 95866 529174
rect 96102 528938 96134 529174
rect 95514 528854 96134 528938
rect 95514 528618 95546 528854
rect 95782 528618 95866 528854
rect 96102 528618 96134 528854
rect 95514 493174 96134 528618
rect 95514 492938 95546 493174
rect 95782 492938 95866 493174
rect 96102 492938 96134 493174
rect 95514 492854 96134 492938
rect 95514 492618 95546 492854
rect 95782 492618 95866 492854
rect 96102 492618 96134 492854
rect 95514 457174 96134 492618
rect 95514 456938 95546 457174
rect 95782 456938 95866 457174
rect 96102 456938 96134 457174
rect 95514 456854 96134 456938
rect 95514 456618 95546 456854
rect 95782 456618 95866 456854
rect 96102 456618 96134 456854
rect 95514 421174 96134 456618
rect 95514 420938 95546 421174
rect 95782 420938 95866 421174
rect 96102 420938 96134 421174
rect 95514 420854 96134 420938
rect 95514 420618 95546 420854
rect 95782 420618 95866 420854
rect 96102 420618 96134 420854
rect 95514 385174 96134 420618
rect 95514 384938 95546 385174
rect 95782 384938 95866 385174
rect 96102 384938 96134 385174
rect 95514 384854 96134 384938
rect 95514 384618 95546 384854
rect 95782 384618 95866 384854
rect 96102 384618 96134 384854
rect 95514 349174 96134 384618
rect 95514 348938 95546 349174
rect 95782 348938 95866 349174
rect 96102 348938 96134 349174
rect 95514 348854 96134 348938
rect 95514 348618 95546 348854
rect 95782 348618 95866 348854
rect 96102 348618 96134 348854
rect 95514 313174 96134 348618
rect 95514 312938 95546 313174
rect 95782 312938 95866 313174
rect 96102 312938 96134 313174
rect 95514 312854 96134 312938
rect 95514 312618 95546 312854
rect 95782 312618 95866 312854
rect 96102 312618 96134 312854
rect 95514 277174 96134 312618
rect 95514 276938 95546 277174
rect 95782 276938 95866 277174
rect 96102 276938 96134 277174
rect 95514 276854 96134 276938
rect 95514 276618 95546 276854
rect 95782 276618 95866 276854
rect 96102 276618 96134 276854
rect 95514 241174 96134 276618
rect 95514 240938 95546 241174
rect 95782 240938 95866 241174
rect 96102 240938 96134 241174
rect 95514 240854 96134 240938
rect 95514 240618 95546 240854
rect 95782 240618 95866 240854
rect 96102 240618 96134 240854
rect 95514 205174 96134 240618
rect 95514 204938 95546 205174
rect 95782 204938 95866 205174
rect 96102 204938 96134 205174
rect 95514 204854 96134 204938
rect 95514 204618 95546 204854
rect 95782 204618 95866 204854
rect 96102 204618 96134 204854
rect 95514 169174 96134 204618
rect 95514 168938 95546 169174
rect 95782 168938 95866 169174
rect 96102 168938 96134 169174
rect 95514 168854 96134 168938
rect 95514 168618 95546 168854
rect 95782 168618 95866 168854
rect 96102 168618 96134 168854
rect 95514 133174 96134 168618
rect 95514 132938 95546 133174
rect 95782 132938 95866 133174
rect 96102 132938 96134 133174
rect 95514 132854 96134 132938
rect 95514 132618 95546 132854
rect 95782 132618 95866 132854
rect 96102 132618 96134 132854
rect 95514 97174 96134 132618
rect 95514 96938 95546 97174
rect 95782 96938 95866 97174
rect 96102 96938 96134 97174
rect 95514 96854 96134 96938
rect 95514 96618 95546 96854
rect 95782 96618 95866 96854
rect 96102 96618 96134 96854
rect 95514 61174 96134 96618
rect 95514 60938 95546 61174
rect 95782 60938 95866 61174
rect 96102 60938 96134 61174
rect 95514 60854 96134 60938
rect 95514 60618 95546 60854
rect 95782 60618 95866 60854
rect 96102 60618 96134 60854
rect 95514 25174 96134 60618
rect 95514 24938 95546 25174
rect 95782 24938 95866 25174
rect 96102 24938 96134 25174
rect 95514 24854 96134 24938
rect 95514 24618 95546 24854
rect 95782 24618 95866 24854
rect 96102 24618 96134 24854
rect 95514 -3226 96134 24618
rect 95514 -3462 95546 -3226
rect 95782 -3462 95866 -3226
rect 96102 -3462 96134 -3226
rect 95514 -3546 96134 -3462
rect 95514 -3782 95546 -3546
rect 95782 -3782 95866 -3546
rect 96102 -3782 96134 -3546
rect 95514 -3814 96134 -3782
rect 99234 676894 99854 709082
rect 99234 676658 99266 676894
rect 99502 676658 99586 676894
rect 99822 676658 99854 676894
rect 99234 676574 99854 676658
rect 99234 676338 99266 676574
rect 99502 676338 99586 676574
rect 99822 676338 99854 676574
rect 99234 640894 99854 676338
rect 99234 640658 99266 640894
rect 99502 640658 99586 640894
rect 99822 640658 99854 640894
rect 99234 640574 99854 640658
rect 99234 640338 99266 640574
rect 99502 640338 99586 640574
rect 99822 640338 99854 640574
rect 99234 604894 99854 640338
rect 99234 604658 99266 604894
rect 99502 604658 99586 604894
rect 99822 604658 99854 604894
rect 99234 604574 99854 604658
rect 99234 604338 99266 604574
rect 99502 604338 99586 604574
rect 99822 604338 99854 604574
rect 99234 568894 99854 604338
rect 99234 568658 99266 568894
rect 99502 568658 99586 568894
rect 99822 568658 99854 568894
rect 99234 568574 99854 568658
rect 99234 568338 99266 568574
rect 99502 568338 99586 568574
rect 99822 568338 99854 568574
rect 99234 532894 99854 568338
rect 99234 532658 99266 532894
rect 99502 532658 99586 532894
rect 99822 532658 99854 532894
rect 99234 532574 99854 532658
rect 99234 532338 99266 532574
rect 99502 532338 99586 532574
rect 99822 532338 99854 532574
rect 99234 496894 99854 532338
rect 99234 496658 99266 496894
rect 99502 496658 99586 496894
rect 99822 496658 99854 496894
rect 99234 496574 99854 496658
rect 99234 496338 99266 496574
rect 99502 496338 99586 496574
rect 99822 496338 99854 496574
rect 99234 460894 99854 496338
rect 99234 460658 99266 460894
rect 99502 460658 99586 460894
rect 99822 460658 99854 460894
rect 99234 460574 99854 460658
rect 99234 460338 99266 460574
rect 99502 460338 99586 460574
rect 99822 460338 99854 460574
rect 99234 424894 99854 460338
rect 99234 424658 99266 424894
rect 99502 424658 99586 424894
rect 99822 424658 99854 424894
rect 99234 424574 99854 424658
rect 99234 424338 99266 424574
rect 99502 424338 99586 424574
rect 99822 424338 99854 424574
rect 99234 388894 99854 424338
rect 99234 388658 99266 388894
rect 99502 388658 99586 388894
rect 99822 388658 99854 388894
rect 99234 388574 99854 388658
rect 99234 388338 99266 388574
rect 99502 388338 99586 388574
rect 99822 388338 99854 388574
rect 99234 352894 99854 388338
rect 99234 352658 99266 352894
rect 99502 352658 99586 352894
rect 99822 352658 99854 352894
rect 99234 352574 99854 352658
rect 99234 352338 99266 352574
rect 99502 352338 99586 352574
rect 99822 352338 99854 352574
rect 99234 316894 99854 352338
rect 99234 316658 99266 316894
rect 99502 316658 99586 316894
rect 99822 316658 99854 316894
rect 99234 316574 99854 316658
rect 99234 316338 99266 316574
rect 99502 316338 99586 316574
rect 99822 316338 99854 316574
rect 99234 280894 99854 316338
rect 99234 280658 99266 280894
rect 99502 280658 99586 280894
rect 99822 280658 99854 280894
rect 99234 280574 99854 280658
rect 99234 280338 99266 280574
rect 99502 280338 99586 280574
rect 99822 280338 99854 280574
rect 99234 244894 99854 280338
rect 99234 244658 99266 244894
rect 99502 244658 99586 244894
rect 99822 244658 99854 244894
rect 99234 244574 99854 244658
rect 99234 244338 99266 244574
rect 99502 244338 99586 244574
rect 99822 244338 99854 244574
rect 99234 208894 99854 244338
rect 99234 208658 99266 208894
rect 99502 208658 99586 208894
rect 99822 208658 99854 208894
rect 99234 208574 99854 208658
rect 99234 208338 99266 208574
rect 99502 208338 99586 208574
rect 99822 208338 99854 208574
rect 99234 172894 99854 208338
rect 99234 172658 99266 172894
rect 99502 172658 99586 172894
rect 99822 172658 99854 172894
rect 99234 172574 99854 172658
rect 99234 172338 99266 172574
rect 99502 172338 99586 172574
rect 99822 172338 99854 172574
rect 99234 136894 99854 172338
rect 99234 136658 99266 136894
rect 99502 136658 99586 136894
rect 99822 136658 99854 136894
rect 99234 136574 99854 136658
rect 99234 136338 99266 136574
rect 99502 136338 99586 136574
rect 99822 136338 99854 136574
rect 99234 100894 99854 136338
rect 99234 100658 99266 100894
rect 99502 100658 99586 100894
rect 99822 100658 99854 100894
rect 99234 100574 99854 100658
rect 99234 100338 99266 100574
rect 99502 100338 99586 100574
rect 99822 100338 99854 100574
rect 99234 64894 99854 100338
rect 99234 64658 99266 64894
rect 99502 64658 99586 64894
rect 99822 64658 99854 64894
rect 99234 64574 99854 64658
rect 99234 64338 99266 64574
rect 99502 64338 99586 64574
rect 99822 64338 99854 64574
rect 99234 28894 99854 64338
rect 99234 28658 99266 28894
rect 99502 28658 99586 28894
rect 99822 28658 99854 28894
rect 99234 28574 99854 28658
rect 99234 28338 99266 28574
rect 99502 28338 99586 28574
rect 99822 28338 99854 28574
rect 99234 -5146 99854 28338
rect 99234 -5382 99266 -5146
rect 99502 -5382 99586 -5146
rect 99822 -5382 99854 -5146
rect 99234 -5466 99854 -5382
rect 99234 -5702 99266 -5466
rect 99502 -5702 99586 -5466
rect 99822 -5702 99854 -5466
rect 99234 -5734 99854 -5702
rect 102954 680614 103574 711002
rect 120954 710598 121574 711590
rect 120954 710362 120986 710598
rect 121222 710362 121306 710598
rect 121542 710362 121574 710598
rect 120954 710278 121574 710362
rect 120954 710042 120986 710278
rect 121222 710042 121306 710278
rect 121542 710042 121574 710278
rect 117234 708678 117854 709670
rect 117234 708442 117266 708678
rect 117502 708442 117586 708678
rect 117822 708442 117854 708678
rect 117234 708358 117854 708442
rect 117234 708122 117266 708358
rect 117502 708122 117586 708358
rect 117822 708122 117854 708358
rect 113514 706758 114134 707750
rect 113514 706522 113546 706758
rect 113782 706522 113866 706758
rect 114102 706522 114134 706758
rect 113514 706438 114134 706522
rect 113514 706202 113546 706438
rect 113782 706202 113866 706438
rect 114102 706202 114134 706438
rect 102954 680378 102986 680614
rect 103222 680378 103306 680614
rect 103542 680378 103574 680614
rect 102954 680294 103574 680378
rect 102954 680058 102986 680294
rect 103222 680058 103306 680294
rect 103542 680058 103574 680294
rect 102954 644614 103574 680058
rect 102954 644378 102986 644614
rect 103222 644378 103306 644614
rect 103542 644378 103574 644614
rect 102954 644294 103574 644378
rect 102954 644058 102986 644294
rect 103222 644058 103306 644294
rect 103542 644058 103574 644294
rect 102954 608614 103574 644058
rect 102954 608378 102986 608614
rect 103222 608378 103306 608614
rect 103542 608378 103574 608614
rect 102954 608294 103574 608378
rect 102954 608058 102986 608294
rect 103222 608058 103306 608294
rect 103542 608058 103574 608294
rect 102954 572614 103574 608058
rect 102954 572378 102986 572614
rect 103222 572378 103306 572614
rect 103542 572378 103574 572614
rect 102954 572294 103574 572378
rect 102954 572058 102986 572294
rect 103222 572058 103306 572294
rect 103542 572058 103574 572294
rect 102954 536614 103574 572058
rect 102954 536378 102986 536614
rect 103222 536378 103306 536614
rect 103542 536378 103574 536614
rect 102954 536294 103574 536378
rect 102954 536058 102986 536294
rect 103222 536058 103306 536294
rect 103542 536058 103574 536294
rect 102954 500614 103574 536058
rect 102954 500378 102986 500614
rect 103222 500378 103306 500614
rect 103542 500378 103574 500614
rect 102954 500294 103574 500378
rect 102954 500058 102986 500294
rect 103222 500058 103306 500294
rect 103542 500058 103574 500294
rect 102954 464614 103574 500058
rect 102954 464378 102986 464614
rect 103222 464378 103306 464614
rect 103542 464378 103574 464614
rect 102954 464294 103574 464378
rect 102954 464058 102986 464294
rect 103222 464058 103306 464294
rect 103542 464058 103574 464294
rect 102954 428614 103574 464058
rect 102954 428378 102986 428614
rect 103222 428378 103306 428614
rect 103542 428378 103574 428614
rect 102954 428294 103574 428378
rect 102954 428058 102986 428294
rect 103222 428058 103306 428294
rect 103542 428058 103574 428294
rect 102954 392614 103574 428058
rect 102954 392378 102986 392614
rect 103222 392378 103306 392614
rect 103542 392378 103574 392614
rect 102954 392294 103574 392378
rect 102954 392058 102986 392294
rect 103222 392058 103306 392294
rect 103542 392058 103574 392294
rect 102954 356614 103574 392058
rect 102954 356378 102986 356614
rect 103222 356378 103306 356614
rect 103542 356378 103574 356614
rect 102954 356294 103574 356378
rect 102954 356058 102986 356294
rect 103222 356058 103306 356294
rect 103542 356058 103574 356294
rect 102954 320614 103574 356058
rect 102954 320378 102986 320614
rect 103222 320378 103306 320614
rect 103542 320378 103574 320614
rect 102954 320294 103574 320378
rect 102954 320058 102986 320294
rect 103222 320058 103306 320294
rect 103542 320058 103574 320294
rect 102954 284614 103574 320058
rect 102954 284378 102986 284614
rect 103222 284378 103306 284614
rect 103542 284378 103574 284614
rect 102954 284294 103574 284378
rect 102954 284058 102986 284294
rect 103222 284058 103306 284294
rect 103542 284058 103574 284294
rect 102954 248614 103574 284058
rect 102954 248378 102986 248614
rect 103222 248378 103306 248614
rect 103542 248378 103574 248614
rect 102954 248294 103574 248378
rect 102954 248058 102986 248294
rect 103222 248058 103306 248294
rect 103542 248058 103574 248294
rect 102954 212614 103574 248058
rect 102954 212378 102986 212614
rect 103222 212378 103306 212614
rect 103542 212378 103574 212614
rect 102954 212294 103574 212378
rect 102954 212058 102986 212294
rect 103222 212058 103306 212294
rect 103542 212058 103574 212294
rect 102954 176614 103574 212058
rect 102954 176378 102986 176614
rect 103222 176378 103306 176614
rect 103542 176378 103574 176614
rect 102954 176294 103574 176378
rect 102954 176058 102986 176294
rect 103222 176058 103306 176294
rect 103542 176058 103574 176294
rect 102954 140614 103574 176058
rect 102954 140378 102986 140614
rect 103222 140378 103306 140614
rect 103542 140378 103574 140614
rect 102954 140294 103574 140378
rect 102954 140058 102986 140294
rect 103222 140058 103306 140294
rect 103542 140058 103574 140294
rect 102954 104614 103574 140058
rect 102954 104378 102986 104614
rect 103222 104378 103306 104614
rect 103542 104378 103574 104614
rect 102954 104294 103574 104378
rect 102954 104058 102986 104294
rect 103222 104058 103306 104294
rect 103542 104058 103574 104294
rect 102954 68614 103574 104058
rect 102954 68378 102986 68614
rect 103222 68378 103306 68614
rect 103542 68378 103574 68614
rect 102954 68294 103574 68378
rect 102954 68058 102986 68294
rect 103222 68058 103306 68294
rect 103542 68058 103574 68294
rect 102954 32614 103574 68058
rect 102954 32378 102986 32614
rect 103222 32378 103306 32614
rect 103542 32378 103574 32614
rect 102954 32294 103574 32378
rect 102954 32058 102986 32294
rect 103222 32058 103306 32294
rect 103542 32058 103574 32294
rect 84954 -6342 84986 -6106
rect 85222 -6342 85306 -6106
rect 85542 -6342 85574 -6106
rect 84954 -6426 85574 -6342
rect 84954 -6662 84986 -6426
rect 85222 -6662 85306 -6426
rect 85542 -6662 85574 -6426
rect 84954 -7654 85574 -6662
rect 102954 -7066 103574 32058
rect 109794 704838 110414 705830
rect 109794 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 110414 704838
rect 109794 704518 110414 704602
rect 109794 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 110414 704518
rect 109794 687454 110414 704282
rect 109794 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 110414 687454
rect 109794 687134 110414 687218
rect 109794 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 110414 687134
rect 109794 651454 110414 686898
rect 109794 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 110414 651454
rect 109794 651134 110414 651218
rect 109794 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 110414 651134
rect 109794 615454 110414 650898
rect 109794 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 110414 615454
rect 109794 615134 110414 615218
rect 109794 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 110414 615134
rect 109794 579454 110414 614898
rect 109794 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 110414 579454
rect 109794 579134 110414 579218
rect 109794 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 110414 579134
rect 109794 543454 110414 578898
rect 109794 543218 109826 543454
rect 110062 543218 110146 543454
rect 110382 543218 110414 543454
rect 109794 543134 110414 543218
rect 109794 542898 109826 543134
rect 110062 542898 110146 543134
rect 110382 542898 110414 543134
rect 109794 507454 110414 542898
rect 109794 507218 109826 507454
rect 110062 507218 110146 507454
rect 110382 507218 110414 507454
rect 109794 507134 110414 507218
rect 109794 506898 109826 507134
rect 110062 506898 110146 507134
rect 110382 506898 110414 507134
rect 109794 471454 110414 506898
rect 109794 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 110414 471454
rect 109794 471134 110414 471218
rect 109794 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 110414 471134
rect 109794 435454 110414 470898
rect 109794 435218 109826 435454
rect 110062 435218 110146 435454
rect 110382 435218 110414 435454
rect 109794 435134 110414 435218
rect 109794 434898 109826 435134
rect 110062 434898 110146 435134
rect 110382 434898 110414 435134
rect 109794 399454 110414 434898
rect 109794 399218 109826 399454
rect 110062 399218 110146 399454
rect 110382 399218 110414 399454
rect 109794 399134 110414 399218
rect 109794 398898 109826 399134
rect 110062 398898 110146 399134
rect 110382 398898 110414 399134
rect 109794 363454 110414 398898
rect 109794 363218 109826 363454
rect 110062 363218 110146 363454
rect 110382 363218 110414 363454
rect 109794 363134 110414 363218
rect 109794 362898 109826 363134
rect 110062 362898 110146 363134
rect 110382 362898 110414 363134
rect 109794 327454 110414 362898
rect 109794 327218 109826 327454
rect 110062 327218 110146 327454
rect 110382 327218 110414 327454
rect 109794 327134 110414 327218
rect 109794 326898 109826 327134
rect 110062 326898 110146 327134
rect 110382 326898 110414 327134
rect 109794 291454 110414 326898
rect 109794 291218 109826 291454
rect 110062 291218 110146 291454
rect 110382 291218 110414 291454
rect 109794 291134 110414 291218
rect 109794 290898 109826 291134
rect 110062 290898 110146 291134
rect 110382 290898 110414 291134
rect 109794 255454 110414 290898
rect 109794 255218 109826 255454
rect 110062 255218 110146 255454
rect 110382 255218 110414 255454
rect 109794 255134 110414 255218
rect 109794 254898 109826 255134
rect 110062 254898 110146 255134
rect 110382 254898 110414 255134
rect 109794 219454 110414 254898
rect 109794 219218 109826 219454
rect 110062 219218 110146 219454
rect 110382 219218 110414 219454
rect 109794 219134 110414 219218
rect 109794 218898 109826 219134
rect 110062 218898 110146 219134
rect 110382 218898 110414 219134
rect 109794 183454 110414 218898
rect 109794 183218 109826 183454
rect 110062 183218 110146 183454
rect 110382 183218 110414 183454
rect 109794 183134 110414 183218
rect 109794 182898 109826 183134
rect 110062 182898 110146 183134
rect 110382 182898 110414 183134
rect 109794 147454 110414 182898
rect 109794 147218 109826 147454
rect 110062 147218 110146 147454
rect 110382 147218 110414 147454
rect 109794 147134 110414 147218
rect 109794 146898 109826 147134
rect 110062 146898 110146 147134
rect 110382 146898 110414 147134
rect 109794 111454 110414 146898
rect 109794 111218 109826 111454
rect 110062 111218 110146 111454
rect 110382 111218 110414 111454
rect 109794 111134 110414 111218
rect 109794 110898 109826 111134
rect 110062 110898 110146 111134
rect 110382 110898 110414 111134
rect 109794 75454 110414 110898
rect 109794 75218 109826 75454
rect 110062 75218 110146 75454
rect 110382 75218 110414 75454
rect 109794 75134 110414 75218
rect 109794 74898 109826 75134
rect 110062 74898 110146 75134
rect 110382 74898 110414 75134
rect 109794 39454 110414 74898
rect 109794 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 110414 39454
rect 109794 39134 110414 39218
rect 109794 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 110414 39134
rect 109794 3454 110414 38898
rect 109794 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 110414 3454
rect 109794 3134 110414 3218
rect 109794 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 110414 3134
rect 109794 -346 110414 2898
rect 109794 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 110414 -346
rect 109794 -666 110414 -582
rect 109794 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 110414 -666
rect 109794 -1894 110414 -902
rect 113514 691174 114134 706202
rect 113514 690938 113546 691174
rect 113782 690938 113866 691174
rect 114102 690938 114134 691174
rect 113514 690854 114134 690938
rect 113514 690618 113546 690854
rect 113782 690618 113866 690854
rect 114102 690618 114134 690854
rect 113514 655174 114134 690618
rect 113514 654938 113546 655174
rect 113782 654938 113866 655174
rect 114102 654938 114134 655174
rect 113514 654854 114134 654938
rect 113514 654618 113546 654854
rect 113782 654618 113866 654854
rect 114102 654618 114134 654854
rect 113514 619174 114134 654618
rect 113514 618938 113546 619174
rect 113782 618938 113866 619174
rect 114102 618938 114134 619174
rect 113514 618854 114134 618938
rect 113514 618618 113546 618854
rect 113782 618618 113866 618854
rect 114102 618618 114134 618854
rect 113514 583174 114134 618618
rect 113514 582938 113546 583174
rect 113782 582938 113866 583174
rect 114102 582938 114134 583174
rect 113514 582854 114134 582938
rect 113514 582618 113546 582854
rect 113782 582618 113866 582854
rect 114102 582618 114134 582854
rect 113514 547174 114134 582618
rect 113514 546938 113546 547174
rect 113782 546938 113866 547174
rect 114102 546938 114134 547174
rect 113514 546854 114134 546938
rect 113514 546618 113546 546854
rect 113782 546618 113866 546854
rect 114102 546618 114134 546854
rect 113514 511174 114134 546618
rect 113514 510938 113546 511174
rect 113782 510938 113866 511174
rect 114102 510938 114134 511174
rect 113514 510854 114134 510938
rect 113514 510618 113546 510854
rect 113782 510618 113866 510854
rect 114102 510618 114134 510854
rect 113514 475174 114134 510618
rect 113514 474938 113546 475174
rect 113782 474938 113866 475174
rect 114102 474938 114134 475174
rect 113514 474854 114134 474938
rect 113514 474618 113546 474854
rect 113782 474618 113866 474854
rect 114102 474618 114134 474854
rect 113514 439174 114134 474618
rect 113514 438938 113546 439174
rect 113782 438938 113866 439174
rect 114102 438938 114134 439174
rect 113514 438854 114134 438938
rect 113514 438618 113546 438854
rect 113782 438618 113866 438854
rect 114102 438618 114134 438854
rect 113514 403174 114134 438618
rect 113514 402938 113546 403174
rect 113782 402938 113866 403174
rect 114102 402938 114134 403174
rect 113514 402854 114134 402938
rect 113514 402618 113546 402854
rect 113782 402618 113866 402854
rect 114102 402618 114134 402854
rect 113514 367174 114134 402618
rect 113514 366938 113546 367174
rect 113782 366938 113866 367174
rect 114102 366938 114134 367174
rect 113514 366854 114134 366938
rect 113514 366618 113546 366854
rect 113782 366618 113866 366854
rect 114102 366618 114134 366854
rect 113514 331174 114134 366618
rect 113514 330938 113546 331174
rect 113782 330938 113866 331174
rect 114102 330938 114134 331174
rect 113514 330854 114134 330938
rect 113514 330618 113546 330854
rect 113782 330618 113866 330854
rect 114102 330618 114134 330854
rect 113514 295174 114134 330618
rect 113514 294938 113546 295174
rect 113782 294938 113866 295174
rect 114102 294938 114134 295174
rect 113514 294854 114134 294938
rect 113514 294618 113546 294854
rect 113782 294618 113866 294854
rect 114102 294618 114134 294854
rect 113514 259174 114134 294618
rect 113514 258938 113546 259174
rect 113782 258938 113866 259174
rect 114102 258938 114134 259174
rect 113514 258854 114134 258938
rect 113514 258618 113546 258854
rect 113782 258618 113866 258854
rect 114102 258618 114134 258854
rect 113514 223174 114134 258618
rect 113514 222938 113546 223174
rect 113782 222938 113866 223174
rect 114102 222938 114134 223174
rect 113514 222854 114134 222938
rect 113514 222618 113546 222854
rect 113782 222618 113866 222854
rect 114102 222618 114134 222854
rect 113514 187174 114134 222618
rect 113514 186938 113546 187174
rect 113782 186938 113866 187174
rect 114102 186938 114134 187174
rect 113514 186854 114134 186938
rect 113514 186618 113546 186854
rect 113782 186618 113866 186854
rect 114102 186618 114134 186854
rect 113514 151174 114134 186618
rect 113514 150938 113546 151174
rect 113782 150938 113866 151174
rect 114102 150938 114134 151174
rect 113514 150854 114134 150938
rect 113514 150618 113546 150854
rect 113782 150618 113866 150854
rect 114102 150618 114134 150854
rect 113514 115174 114134 150618
rect 113514 114938 113546 115174
rect 113782 114938 113866 115174
rect 114102 114938 114134 115174
rect 113514 114854 114134 114938
rect 113514 114618 113546 114854
rect 113782 114618 113866 114854
rect 114102 114618 114134 114854
rect 113514 79174 114134 114618
rect 113514 78938 113546 79174
rect 113782 78938 113866 79174
rect 114102 78938 114134 79174
rect 113514 78854 114134 78938
rect 113514 78618 113546 78854
rect 113782 78618 113866 78854
rect 114102 78618 114134 78854
rect 113514 43174 114134 78618
rect 113514 42938 113546 43174
rect 113782 42938 113866 43174
rect 114102 42938 114134 43174
rect 113514 42854 114134 42938
rect 113514 42618 113546 42854
rect 113782 42618 113866 42854
rect 114102 42618 114134 42854
rect 113514 7174 114134 42618
rect 113514 6938 113546 7174
rect 113782 6938 113866 7174
rect 114102 6938 114134 7174
rect 113514 6854 114134 6938
rect 113514 6618 113546 6854
rect 113782 6618 113866 6854
rect 114102 6618 114134 6854
rect 113514 -2266 114134 6618
rect 113514 -2502 113546 -2266
rect 113782 -2502 113866 -2266
rect 114102 -2502 114134 -2266
rect 113514 -2586 114134 -2502
rect 113514 -2822 113546 -2586
rect 113782 -2822 113866 -2586
rect 114102 -2822 114134 -2586
rect 113514 -3814 114134 -2822
rect 117234 694894 117854 708122
rect 117234 694658 117266 694894
rect 117502 694658 117586 694894
rect 117822 694658 117854 694894
rect 117234 694574 117854 694658
rect 117234 694338 117266 694574
rect 117502 694338 117586 694574
rect 117822 694338 117854 694574
rect 117234 658894 117854 694338
rect 117234 658658 117266 658894
rect 117502 658658 117586 658894
rect 117822 658658 117854 658894
rect 117234 658574 117854 658658
rect 117234 658338 117266 658574
rect 117502 658338 117586 658574
rect 117822 658338 117854 658574
rect 117234 622894 117854 658338
rect 117234 622658 117266 622894
rect 117502 622658 117586 622894
rect 117822 622658 117854 622894
rect 117234 622574 117854 622658
rect 117234 622338 117266 622574
rect 117502 622338 117586 622574
rect 117822 622338 117854 622574
rect 117234 586894 117854 622338
rect 117234 586658 117266 586894
rect 117502 586658 117586 586894
rect 117822 586658 117854 586894
rect 117234 586574 117854 586658
rect 117234 586338 117266 586574
rect 117502 586338 117586 586574
rect 117822 586338 117854 586574
rect 117234 550894 117854 586338
rect 117234 550658 117266 550894
rect 117502 550658 117586 550894
rect 117822 550658 117854 550894
rect 117234 550574 117854 550658
rect 117234 550338 117266 550574
rect 117502 550338 117586 550574
rect 117822 550338 117854 550574
rect 117234 514894 117854 550338
rect 117234 514658 117266 514894
rect 117502 514658 117586 514894
rect 117822 514658 117854 514894
rect 117234 514574 117854 514658
rect 117234 514338 117266 514574
rect 117502 514338 117586 514574
rect 117822 514338 117854 514574
rect 117234 478894 117854 514338
rect 117234 478658 117266 478894
rect 117502 478658 117586 478894
rect 117822 478658 117854 478894
rect 117234 478574 117854 478658
rect 117234 478338 117266 478574
rect 117502 478338 117586 478574
rect 117822 478338 117854 478574
rect 117234 442894 117854 478338
rect 117234 442658 117266 442894
rect 117502 442658 117586 442894
rect 117822 442658 117854 442894
rect 117234 442574 117854 442658
rect 117234 442338 117266 442574
rect 117502 442338 117586 442574
rect 117822 442338 117854 442574
rect 117234 406894 117854 442338
rect 117234 406658 117266 406894
rect 117502 406658 117586 406894
rect 117822 406658 117854 406894
rect 117234 406574 117854 406658
rect 117234 406338 117266 406574
rect 117502 406338 117586 406574
rect 117822 406338 117854 406574
rect 117234 370894 117854 406338
rect 117234 370658 117266 370894
rect 117502 370658 117586 370894
rect 117822 370658 117854 370894
rect 117234 370574 117854 370658
rect 117234 370338 117266 370574
rect 117502 370338 117586 370574
rect 117822 370338 117854 370574
rect 117234 334894 117854 370338
rect 117234 334658 117266 334894
rect 117502 334658 117586 334894
rect 117822 334658 117854 334894
rect 117234 334574 117854 334658
rect 117234 334338 117266 334574
rect 117502 334338 117586 334574
rect 117822 334338 117854 334574
rect 117234 298894 117854 334338
rect 117234 298658 117266 298894
rect 117502 298658 117586 298894
rect 117822 298658 117854 298894
rect 117234 298574 117854 298658
rect 117234 298338 117266 298574
rect 117502 298338 117586 298574
rect 117822 298338 117854 298574
rect 117234 262894 117854 298338
rect 117234 262658 117266 262894
rect 117502 262658 117586 262894
rect 117822 262658 117854 262894
rect 117234 262574 117854 262658
rect 117234 262338 117266 262574
rect 117502 262338 117586 262574
rect 117822 262338 117854 262574
rect 117234 226894 117854 262338
rect 117234 226658 117266 226894
rect 117502 226658 117586 226894
rect 117822 226658 117854 226894
rect 117234 226574 117854 226658
rect 117234 226338 117266 226574
rect 117502 226338 117586 226574
rect 117822 226338 117854 226574
rect 117234 190894 117854 226338
rect 117234 190658 117266 190894
rect 117502 190658 117586 190894
rect 117822 190658 117854 190894
rect 117234 190574 117854 190658
rect 117234 190338 117266 190574
rect 117502 190338 117586 190574
rect 117822 190338 117854 190574
rect 117234 154894 117854 190338
rect 117234 154658 117266 154894
rect 117502 154658 117586 154894
rect 117822 154658 117854 154894
rect 117234 154574 117854 154658
rect 117234 154338 117266 154574
rect 117502 154338 117586 154574
rect 117822 154338 117854 154574
rect 117234 118894 117854 154338
rect 117234 118658 117266 118894
rect 117502 118658 117586 118894
rect 117822 118658 117854 118894
rect 117234 118574 117854 118658
rect 117234 118338 117266 118574
rect 117502 118338 117586 118574
rect 117822 118338 117854 118574
rect 117234 82894 117854 118338
rect 117234 82658 117266 82894
rect 117502 82658 117586 82894
rect 117822 82658 117854 82894
rect 117234 82574 117854 82658
rect 117234 82338 117266 82574
rect 117502 82338 117586 82574
rect 117822 82338 117854 82574
rect 117234 46894 117854 82338
rect 117234 46658 117266 46894
rect 117502 46658 117586 46894
rect 117822 46658 117854 46894
rect 117234 46574 117854 46658
rect 117234 46338 117266 46574
rect 117502 46338 117586 46574
rect 117822 46338 117854 46574
rect 117234 10894 117854 46338
rect 117234 10658 117266 10894
rect 117502 10658 117586 10894
rect 117822 10658 117854 10894
rect 117234 10574 117854 10658
rect 117234 10338 117266 10574
rect 117502 10338 117586 10574
rect 117822 10338 117854 10574
rect 117234 -4186 117854 10338
rect 117234 -4422 117266 -4186
rect 117502 -4422 117586 -4186
rect 117822 -4422 117854 -4186
rect 117234 -4506 117854 -4422
rect 117234 -4742 117266 -4506
rect 117502 -4742 117586 -4506
rect 117822 -4742 117854 -4506
rect 117234 -5734 117854 -4742
rect 120954 698614 121574 710042
rect 138954 711558 139574 711590
rect 138954 711322 138986 711558
rect 139222 711322 139306 711558
rect 139542 711322 139574 711558
rect 138954 711238 139574 711322
rect 138954 711002 138986 711238
rect 139222 711002 139306 711238
rect 139542 711002 139574 711238
rect 135234 709638 135854 709670
rect 135234 709402 135266 709638
rect 135502 709402 135586 709638
rect 135822 709402 135854 709638
rect 135234 709318 135854 709402
rect 135234 709082 135266 709318
rect 135502 709082 135586 709318
rect 135822 709082 135854 709318
rect 131514 707718 132134 707750
rect 131514 707482 131546 707718
rect 131782 707482 131866 707718
rect 132102 707482 132134 707718
rect 131514 707398 132134 707482
rect 131514 707162 131546 707398
rect 131782 707162 131866 707398
rect 132102 707162 132134 707398
rect 120954 698378 120986 698614
rect 121222 698378 121306 698614
rect 121542 698378 121574 698614
rect 120954 698294 121574 698378
rect 120954 698058 120986 698294
rect 121222 698058 121306 698294
rect 121542 698058 121574 698294
rect 120954 662614 121574 698058
rect 120954 662378 120986 662614
rect 121222 662378 121306 662614
rect 121542 662378 121574 662614
rect 120954 662294 121574 662378
rect 120954 662058 120986 662294
rect 121222 662058 121306 662294
rect 121542 662058 121574 662294
rect 120954 626614 121574 662058
rect 120954 626378 120986 626614
rect 121222 626378 121306 626614
rect 121542 626378 121574 626614
rect 120954 626294 121574 626378
rect 120954 626058 120986 626294
rect 121222 626058 121306 626294
rect 121542 626058 121574 626294
rect 120954 590614 121574 626058
rect 120954 590378 120986 590614
rect 121222 590378 121306 590614
rect 121542 590378 121574 590614
rect 120954 590294 121574 590378
rect 120954 590058 120986 590294
rect 121222 590058 121306 590294
rect 121542 590058 121574 590294
rect 120954 554614 121574 590058
rect 120954 554378 120986 554614
rect 121222 554378 121306 554614
rect 121542 554378 121574 554614
rect 120954 554294 121574 554378
rect 120954 554058 120986 554294
rect 121222 554058 121306 554294
rect 121542 554058 121574 554294
rect 120954 518614 121574 554058
rect 120954 518378 120986 518614
rect 121222 518378 121306 518614
rect 121542 518378 121574 518614
rect 120954 518294 121574 518378
rect 120954 518058 120986 518294
rect 121222 518058 121306 518294
rect 121542 518058 121574 518294
rect 120954 482614 121574 518058
rect 120954 482378 120986 482614
rect 121222 482378 121306 482614
rect 121542 482378 121574 482614
rect 120954 482294 121574 482378
rect 120954 482058 120986 482294
rect 121222 482058 121306 482294
rect 121542 482058 121574 482294
rect 120954 446614 121574 482058
rect 120954 446378 120986 446614
rect 121222 446378 121306 446614
rect 121542 446378 121574 446614
rect 120954 446294 121574 446378
rect 120954 446058 120986 446294
rect 121222 446058 121306 446294
rect 121542 446058 121574 446294
rect 120954 410614 121574 446058
rect 120954 410378 120986 410614
rect 121222 410378 121306 410614
rect 121542 410378 121574 410614
rect 120954 410294 121574 410378
rect 120954 410058 120986 410294
rect 121222 410058 121306 410294
rect 121542 410058 121574 410294
rect 120954 374614 121574 410058
rect 120954 374378 120986 374614
rect 121222 374378 121306 374614
rect 121542 374378 121574 374614
rect 120954 374294 121574 374378
rect 120954 374058 120986 374294
rect 121222 374058 121306 374294
rect 121542 374058 121574 374294
rect 120954 338614 121574 374058
rect 120954 338378 120986 338614
rect 121222 338378 121306 338614
rect 121542 338378 121574 338614
rect 120954 338294 121574 338378
rect 120954 338058 120986 338294
rect 121222 338058 121306 338294
rect 121542 338058 121574 338294
rect 120954 302614 121574 338058
rect 120954 302378 120986 302614
rect 121222 302378 121306 302614
rect 121542 302378 121574 302614
rect 120954 302294 121574 302378
rect 120954 302058 120986 302294
rect 121222 302058 121306 302294
rect 121542 302058 121574 302294
rect 120954 266614 121574 302058
rect 120954 266378 120986 266614
rect 121222 266378 121306 266614
rect 121542 266378 121574 266614
rect 120954 266294 121574 266378
rect 120954 266058 120986 266294
rect 121222 266058 121306 266294
rect 121542 266058 121574 266294
rect 120954 230614 121574 266058
rect 120954 230378 120986 230614
rect 121222 230378 121306 230614
rect 121542 230378 121574 230614
rect 120954 230294 121574 230378
rect 120954 230058 120986 230294
rect 121222 230058 121306 230294
rect 121542 230058 121574 230294
rect 120954 194614 121574 230058
rect 120954 194378 120986 194614
rect 121222 194378 121306 194614
rect 121542 194378 121574 194614
rect 120954 194294 121574 194378
rect 120954 194058 120986 194294
rect 121222 194058 121306 194294
rect 121542 194058 121574 194294
rect 120954 158614 121574 194058
rect 120954 158378 120986 158614
rect 121222 158378 121306 158614
rect 121542 158378 121574 158614
rect 120954 158294 121574 158378
rect 120954 158058 120986 158294
rect 121222 158058 121306 158294
rect 121542 158058 121574 158294
rect 120954 122614 121574 158058
rect 120954 122378 120986 122614
rect 121222 122378 121306 122614
rect 121542 122378 121574 122614
rect 120954 122294 121574 122378
rect 120954 122058 120986 122294
rect 121222 122058 121306 122294
rect 121542 122058 121574 122294
rect 120954 86614 121574 122058
rect 120954 86378 120986 86614
rect 121222 86378 121306 86614
rect 121542 86378 121574 86614
rect 120954 86294 121574 86378
rect 120954 86058 120986 86294
rect 121222 86058 121306 86294
rect 121542 86058 121574 86294
rect 120954 50614 121574 86058
rect 120954 50378 120986 50614
rect 121222 50378 121306 50614
rect 121542 50378 121574 50614
rect 120954 50294 121574 50378
rect 120954 50058 120986 50294
rect 121222 50058 121306 50294
rect 121542 50058 121574 50294
rect 120954 14614 121574 50058
rect 120954 14378 120986 14614
rect 121222 14378 121306 14614
rect 121542 14378 121574 14614
rect 120954 14294 121574 14378
rect 120954 14058 120986 14294
rect 121222 14058 121306 14294
rect 121542 14058 121574 14294
rect 102954 -7302 102986 -7066
rect 103222 -7302 103306 -7066
rect 103542 -7302 103574 -7066
rect 102954 -7386 103574 -7302
rect 102954 -7622 102986 -7386
rect 103222 -7622 103306 -7386
rect 103542 -7622 103574 -7386
rect 102954 -7654 103574 -7622
rect 120954 -6106 121574 14058
rect 127794 705798 128414 705830
rect 127794 705562 127826 705798
rect 128062 705562 128146 705798
rect 128382 705562 128414 705798
rect 127794 705478 128414 705562
rect 127794 705242 127826 705478
rect 128062 705242 128146 705478
rect 128382 705242 128414 705478
rect 127794 669454 128414 705242
rect 127794 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 128414 669454
rect 127794 669134 128414 669218
rect 127794 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 128414 669134
rect 127794 633454 128414 668898
rect 127794 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 128414 633454
rect 127794 633134 128414 633218
rect 127794 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 128414 633134
rect 127794 597454 128414 632898
rect 127794 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 128414 597454
rect 127794 597134 128414 597218
rect 127794 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 128414 597134
rect 127794 561454 128414 596898
rect 127794 561218 127826 561454
rect 128062 561218 128146 561454
rect 128382 561218 128414 561454
rect 127794 561134 128414 561218
rect 127794 560898 127826 561134
rect 128062 560898 128146 561134
rect 128382 560898 128414 561134
rect 127794 525454 128414 560898
rect 127794 525218 127826 525454
rect 128062 525218 128146 525454
rect 128382 525218 128414 525454
rect 127794 525134 128414 525218
rect 127794 524898 127826 525134
rect 128062 524898 128146 525134
rect 128382 524898 128414 525134
rect 127794 489454 128414 524898
rect 127794 489218 127826 489454
rect 128062 489218 128146 489454
rect 128382 489218 128414 489454
rect 127794 489134 128414 489218
rect 127794 488898 127826 489134
rect 128062 488898 128146 489134
rect 128382 488898 128414 489134
rect 127794 453454 128414 488898
rect 127794 453218 127826 453454
rect 128062 453218 128146 453454
rect 128382 453218 128414 453454
rect 127794 453134 128414 453218
rect 127794 452898 127826 453134
rect 128062 452898 128146 453134
rect 128382 452898 128414 453134
rect 127794 417454 128414 452898
rect 127794 417218 127826 417454
rect 128062 417218 128146 417454
rect 128382 417218 128414 417454
rect 127794 417134 128414 417218
rect 127794 416898 127826 417134
rect 128062 416898 128146 417134
rect 128382 416898 128414 417134
rect 127794 381454 128414 416898
rect 127794 381218 127826 381454
rect 128062 381218 128146 381454
rect 128382 381218 128414 381454
rect 127794 381134 128414 381218
rect 127794 380898 127826 381134
rect 128062 380898 128146 381134
rect 128382 380898 128414 381134
rect 127794 345454 128414 380898
rect 127794 345218 127826 345454
rect 128062 345218 128146 345454
rect 128382 345218 128414 345454
rect 127794 345134 128414 345218
rect 127794 344898 127826 345134
rect 128062 344898 128146 345134
rect 128382 344898 128414 345134
rect 127794 309454 128414 344898
rect 127794 309218 127826 309454
rect 128062 309218 128146 309454
rect 128382 309218 128414 309454
rect 127794 309134 128414 309218
rect 127794 308898 127826 309134
rect 128062 308898 128146 309134
rect 128382 308898 128414 309134
rect 127794 273454 128414 308898
rect 127794 273218 127826 273454
rect 128062 273218 128146 273454
rect 128382 273218 128414 273454
rect 127794 273134 128414 273218
rect 127794 272898 127826 273134
rect 128062 272898 128146 273134
rect 128382 272898 128414 273134
rect 127794 237454 128414 272898
rect 127794 237218 127826 237454
rect 128062 237218 128146 237454
rect 128382 237218 128414 237454
rect 127794 237134 128414 237218
rect 127794 236898 127826 237134
rect 128062 236898 128146 237134
rect 128382 236898 128414 237134
rect 127794 201454 128414 236898
rect 127794 201218 127826 201454
rect 128062 201218 128146 201454
rect 128382 201218 128414 201454
rect 127794 201134 128414 201218
rect 127794 200898 127826 201134
rect 128062 200898 128146 201134
rect 128382 200898 128414 201134
rect 127794 165454 128414 200898
rect 127794 165218 127826 165454
rect 128062 165218 128146 165454
rect 128382 165218 128414 165454
rect 127794 165134 128414 165218
rect 127794 164898 127826 165134
rect 128062 164898 128146 165134
rect 128382 164898 128414 165134
rect 127794 129454 128414 164898
rect 127794 129218 127826 129454
rect 128062 129218 128146 129454
rect 128382 129218 128414 129454
rect 127794 129134 128414 129218
rect 127794 128898 127826 129134
rect 128062 128898 128146 129134
rect 128382 128898 128414 129134
rect 127794 93454 128414 128898
rect 127794 93218 127826 93454
rect 128062 93218 128146 93454
rect 128382 93218 128414 93454
rect 127794 93134 128414 93218
rect 127794 92898 127826 93134
rect 128062 92898 128146 93134
rect 128382 92898 128414 93134
rect 127794 57454 128414 92898
rect 127794 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 128414 57454
rect 127794 57134 128414 57218
rect 127794 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 128414 57134
rect 127794 21454 128414 56898
rect 127794 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 128414 21454
rect 127794 21134 128414 21218
rect 127794 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 128414 21134
rect 127794 -1306 128414 20898
rect 127794 -1542 127826 -1306
rect 128062 -1542 128146 -1306
rect 128382 -1542 128414 -1306
rect 127794 -1626 128414 -1542
rect 127794 -1862 127826 -1626
rect 128062 -1862 128146 -1626
rect 128382 -1862 128414 -1626
rect 127794 -1894 128414 -1862
rect 131514 673174 132134 707162
rect 131514 672938 131546 673174
rect 131782 672938 131866 673174
rect 132102 672938 132134 673174
rect 131514 672854 132134 672938
rect 131514 672618 131546 672854
rect 131782 672618 131866 672854
rect 132102 672618 132134 672854
rect 131514 637174 132134 672618
rect 131514 636938 131546 637174
rect 131782 636938 131866 637174
rect 132102 636938 132134 637174
rect 131514 636854 132134 636938
rect 131514 636618 131546 636854
rect 131782 636618 131866 636854
rect 132102 636618 132134 636854
rect 131514 601174 132134 636618
rect 131514 600938 131546 601174
rect 131782 600938 131866 601174
rect 132102 600938 132134 601174
rect 131514 600854 132134 600938
rect 131514 600618 131546 600854
rect 131782 600618 131866 600854
rect 132102 600618 132134 600854
rect 131514 565174 132134 600618
rect 131514 564938 131546 565174
rect 131782 564938 131866 565174
rect 132102 564938 132134 565174
rect 131514 564854 132134 564938
rect 131514 564618 131546 564854
rect 131782 564618 131866 564854
rect 132102 564618 132134 564854
rect 131514 529174 132134 564618
rect 131514 528938 131546 529174
rect 131782 528938 131866 529174
rect 132102 528938 132134 529174
rect 131514 528854 132134 528938
rect 131514 528618 131546 528854
rect 131782 528618 131866 528854
rect 132102 528618 132134 528854
rect 131514 493174 132134 528618
rect 131514 492938 131546 493174
rect 131782 492938 131866 493174
rect 132102 492938 132134 493174
rect 131514 492854 132134 492938
rect 131514 492618 131546 492854
rect 131782 492618 131866 492854
rect 132102 492618 132134 492854
rect 131514 457174 132134 492618
rect 131514 456938 131546 457174
rect 131782 456938 131866 457174
rect 132102 456938 132134 457174
rect 131514 456854 132134 456938
rect 131514 456618 131546 456854
rect 131782 456618 131866 456854
rect 132102 456618 132134 456854
rect 131514 421174 132134 456618
rect 131514 420938 131546 421174
rect 131782 420938 131866 421174
rect 132102 420938 132134 421174
rect 131514 420854 132134 420938
rect 131514 420618 131546 420854
rect 131782 420618 131866 420854
rect 132102 420618 132134 420854
rect 131514 385174 132134 420618
rect 131514 384938 131546 385174
rect 131782 384938 131866 385174
rect 132102 384938 132134 385174
rect 131514 384854 132134 384938
rect 131514 384618 131546 384854
rect 131782 384618 131866 384854
rect 132102 384618 132134 384854
rect 131514 349174 132134 384618
rect 131514 348938 131546 349174
rect 131782 348938 131866 349174
rect 132102 348938 132134 349174
rect 131514 348854 132134 348938
rect 131514 348618 131546 348854
rect 131782 348618 131866 348854
rect 132102 348618 132134 348854
rect 131514 313174 132134 348618
rect 131514 312938 131546 313174
rect 131782 312938 131866 313174
rect 132102 312938 132134 313174
rect 131514 312854 132134 312938
rect 131514 312618 131546 312854
rect 131782 312618 131866 312854
rect 132102 312618 132134 312854
rect 131514 277174 132134 312618
rect 131514 276938 131546 277174
rect 131782 276938 131866 277174
rect 132102 276938 132134 277174
rect 131514 276854 132134 276938
rect 131514 276618 131546 276854
rect 131782 276618 131866 276854
rect 132102 276618 132134 276854
rect 131514 241174 132134 276618
rect 131514 240938 131546 241174
rect 131782 240938 131866 241174
rect 132102 240938 132134 241174
rect 131514 240854 132134 240938
rect 131514 240618 131546 240854
rect 131782 240618 131866 240854
rect 132102 240618 132134 240854
rect 131514 205174 132134 240618
rect 131514 204938 131546 205174
rect 131782 204938 131866 205174
rect 132102 204938 132134 205174
rect 131514 204854 132134 204938
rect 131514 204618 131546 204854
rect 131782 204618 131866 204854
rect 132102 204618 132134 204854
rect 131514 169174 132134 204618
rect 131514 168938 131546 169174
rect 131782 168938 131866 169174
rect 132102 168938 132134 169174
rect 131514 168854 132134 168938
rect 131514 168618 131546 168854
rect 131782 168618 131866 168854
rect 132102 168618 132134 168854
rect 131514 133174 132134 168618
rect 131514 132938 131546 133174
rect 131782 132938 131866 133174
rect 132102 132938 132134 133174
rect 131514 132854 132134 132938
rect 131514 132618 131546 132854
rect 131782 132618 131866 132854
rect 132102 132618 132134 132854
rect 131514 97174 132134 132618
rect 131514 96938 131546 97174
rect 131782 96938 131866 97174
rect 132102 96938 132134 97174
rect 131514 96854 132134 96938
rect 131514 96618 131546 96854
rect 131782 96618 131866 96854
rect 132102 96618 132134 96854
rect 131514 61174 132134 96618
rect 131514 60938 131546 61174
rect 131782 60938 131866 61174
rect 132102 60938 132134 61174
rect 131514 60854 132134 60938
rect 131514 60618 131546 60854
rect 131782 60618 131866 60854
rect 132102 60618 132134 60854
rect 131514 25174 132134 60618
rect 131514 24938 131546 25174
rect 131782 24938 131866 25174
rect 132102 24938 132134 25174
rect 131514 24854 132134 24938
rect 131514 24618 131546 24854
rect 131782 24618 131866 24854
rect 132102 24618 132134 24854
rect 131514 -3226 132134 24618
rect 131514 -3462 131546 -3226
rect 131782 -3462 131866 -3226
rect 132102 -3462 132134 -3226
rect 131514 -3546 132134 -3462
rect 131514 -3782 131546 -3546
rect 131782 -3782 131866 -3546
rect 132102 -3782 132134 -3546
rect 131514 -3814 132134 -3782
rect 135234 676894 135854 709082
rect 135234 676658 135266 676894
rect 135502 676658 135586 676894
rect 135822 676658 135854 676894
rect 135234 676574 135854 676658
rect 135234 676338 135266 676574
rect 135502 676338 135586 676574
rect 135822 676338 135854 676574
rect 135234 640894 135854 676338
rect 135234 640658 135266 640894
rect 135502 640658 135586 640894
rect 135822 640658 135854 640894
rect 135234 640574 135854 640658
rect 135234 640338 135266 640574
rect 135502 640338 135586 640574
rect 135822 640338 135854 640574
rect 135234 604894 135854 640338
rect 135234 604658 135266 604894
rect 135502 604658 135586 604894
rect 135822 604658 135854 604894
rect 135234 604574 135854 604658
rect 135234 604338 135266 604574
rect 135502 604338 135586 604574
rect 135822 604338 135854 604574
rect 135234 568894 135854 604338
rect 135234 568658 135266 568894
rect 135502 568658 135586 568894
rect 135822 568658 135854 568894
rect 135234 568574 135854 568658
rect 135234 568338 135266 568574
rect 135502 568338 135586 568574
rect 135822 568338 135854 568574
rect 135234 532894 135854 568338
rect 135234 532658 135266 532894
rect 135502 532658 135586 532894
rect 135822 532658 135854 532894
rect 135234 532574 135854 532658
rect 135234 532338 135266 532574
rect 135502 532338 135586 532574
rect 135822 532338 135854 532574
rect 135234 496894 135854 532338
rect 135234 496658 135266 496894
rect 135502 496658 135586 496894
rect 135822 496658 135854 496894
rect 135234 496574 135854 496658
rect 135234 496338 135266 496574
rect 135502 496338 135586 496574
rect 135822 496338 135854 496574
rect 135234 460894 135854 496338
rect 135234 460658 135266 460894
rect 135502 460658 135586 460894
rect 135822 460658 135854 460894
rect 135234 460574 135854 460658
rect 135234 460338 135266 460574
rect 135502 460338 135586 460574
rect 135822 460338 135854 460574
rect 135234 424894 135854 460338
rect 135234 424658 135266 424894
rect 135502 424658 135586 424894
rect 135822 424658 135854 424894
rect 135234 424574 135854 424658
rect 135234 424338 135266 424574
rect 135502 424338 135586 424574
rect 135822 424338 135854 424574
rect 135234 388894 135854 424338
rect 135234 388658 135266 388894
rect 135502 388658 135586 388894
rect 135822 388658 135854 388894
rect 135234 388574 135854 388658
rect 135234 388338 135266 388574
rect 135502 388338 135586 388574
rect 135822 388338 135854 388574
rect 135234 352894 135854 388338
rect 135234 352658 135266 352894
rect 135502 352658 135586 352894
rect 135822 352658 135854 352894
rect 135234 352574 135854 352658
rect 135234 352338 135266 352574
rect 135502 352338 135586 352574
rect 135822 352338 135854 352574
rect 135234 316894 135854 352338
rect 135234 316658 135266 316894
rect 135502 316658 135586 316894
rect 135822 316658 135854 316894
rect 135234 316574 135854 316658
rect 135234 316338 135266 316574
rect 135502 316338 135586 316574
rect 135822 316338 135854 316574
rect 135234 280894 135854 316338
rect 135234 280658 135266 280894
rect 135502 280658 135586 280894
rect 135822 280658 135854 280894
rect 135234 280574 135854 280658
rect 135234 280338 135266 280574
rect 135502 280338 135586 280574
rect 135822 280338 135854 280574
rect 135234 244894 135854 280338
rect 135234 244658 135266 244894
rect 135502 244658 135586 244894
rect 135822 244658 135854 244894
rect 135234 244574 135854 244658
rect 135234 244338 135266 244574
rect 135502 244338 135586 244574
rect 135822 244338 135854 244574
rect 135234 208894 135854 244338
rect 135234 208658 135266 208894
rect 135502 208658 135586 208894
rect 135822 208658 135854 208894
rect 135234 208574 135854 208658
rect 135234 208338 135266 208574
rect 135502 208338 135586 208574
rect 135822 208338 135854 208574
rect 135234 172894 135854 208338
rect 135234 172658 135266 172894
rect 135502 172658 135586 172894
rect 135822 172658 135854 172894
rect 135234 172574 135854 172658
rect 135234 172338 135266 172574
rect 135502 172338 135586 172574
rect 135822 172338 135854 172574
rect 135234 136894 135854 172338
rect 135234 136658 135266 136894
rect 135502 136658 135586 136894
rect 135822 136658 135854 136894
rect 135234 136574 135854 136658
rect 135234 136338 135266 136574
rect 135502 136338 135586 136574
rect 135822 136338 135854 136574
rect 135234 100894 135854 136338
rect 135234 100658 135266 100894
rect 135502 100658 135586 100894
rect 135822 100658 135854 100894
rect 135234 100574 135854 100658
rect 135234 100338 135266 100574
rect 135502 100338 135586 100574
rect 135822 100338 135854 100574
rect 135234 64894 135854 100338
rect 135234 64658 135266 64894
rect 135502 64658 135586 64894
rect 135822 64658 135854 64894
rect 135234 64574 135854 64658
rect 135234 64338 135266 64574
rect 135502 64338 135586 64574
rect 135822 64338 135854 64574
rect 135234 28894 135854 64338
rect 135234 28658 135266 28894
rect 135502 28658 135586 28894
rect 135822 28658 135854 28894
rect 135234 28574 135854 28658
rect 135234 28338 135266 28574
rect 135502 28338 135586 28574
rect 135822 28338 135854 28574
rect 135234 -5146 135854 28338
rect 135234 -5382 135266 -5146
rect 135502 -5382 135586 -5146
rect 135822 -5382 135854 -5146
rect 135234 -5466 135854 -5382
rect 135234 -5702 135266 -5466
rect 135502 -5702 135586 -5466
rect 135822 -5702 135854 -5466
rect 135234 -5734 135854 -5702
rect 138954 680614 139574 711002
rect 156954 710598 157574 711590
rect 156954 710362 156986 710598
rect 157222 710362 157306 710598
rect 157542 710362 157574 710598
rect 156954 710278 157574 710362
rect 156954 710042 156986 710278
rect 157222 710042 157306 710278
rect 157542 710042 157574 710278
rect 153234 708678 153854 709670
rect 153234 708442 153266 708678
rect 153502 708442 153586 708678
rect 153822 708442 153854 708678
rect 153234 708358 153854 708442
rect 153234 708122 153266 708358
rect 153502 708122 153586 708358
rect 153822 708122 153854 708358
rect 149514 706758 150134 707750
rect 149514 706522 149546 706758
rect 149782 706522 149866 706758
rect 150102 706522 150134 706758
rect 149514 706438 150134 706522
rect 149514 706202 149546 706438
rect 149782 706202 149866 706438
rect 150102 706202 150134 706438
rect 138954 680378 138986 680614
rect 139222 680378 139306 680614
rect 139542 680378 139574 680614
rect 138954 680294 139574 680378
rect 138954 680058 138986 680294
rect 139222 680058 139306 680294
rect 139542 680058 139574 680294
rect 138954 644614 139574 680058
rect 138954 644378 138986 644614
rect 139222 644378 139306 644614
rect 139542 644378 139574 644614
rect 138954 644294 139574 644378
rect 138954 644058 138986 644294
rect 139222 644058 139306 644294
rect 139542 644058 139574 644294
rect 138954 608614 139574 644058
rect 138954 608378 138986 608614
rect 139222 608378 139306 608614
rect 139542 608378 139574 608614
rect 138954 608294 139574 608378
rect 138954 608058 138986 608294
rect 139222 608058 139306 608294
rect 139542 608058 139574 608294
rect 138954 572614 139574 608058
rect 138954 572378 138986 572614
rect 139222 572378 139306 572614
rect 139542 572378 139574 572614
rect 138954 572294 139574 572378
rect 138954 572058 138986 572294
rect 139222 572058 139306 572294
rect 139542 572058 139574 572294
rect 138954 536614 139574 572058
rect 138954 536378 138986 536614
rect 139222 536378 139306 536614
rect 139542 536378 139574 536614
rect 138954 536294 139574 536378
rect 138954 536058 138986 536294
rect 139222 536058 139306 536294
rect 139542 536058 139574 536294
rect 138954 500614 139574 536058
rect 138954 500378 138986 500614
rect 139222 500378 139306 500614
rect 139542 500378 139574 500614
rect 138954 500294 139574 500378
rect 138954 500058 138986 500294
rect 139222 500058 139306 500294
rect 139542 500058 139574 500294
rect 138954 464614 139574 500058
rect 138954 464378 138986 464614
rect 139222 464378 139306 464614
rect 139542 464378 139574 464614
rect 138954 464294 139574 464378
rect 138954 464058 138986 464294
rect 139222 464058 139306 464294
rect 139542 464058 139574 464294
rect 138954 428614 139574 464058
rect 138954 428378 138986 428614
rect 139222 428378 139306 428614
rect 139542 428378 139574 428614
rect 138954 428294 139574 428378
rect 138954 428058 138986 428294
rect 139222 428058 139306 428294
rect 139542 428058 139574 428294
rect 138954 392614 139574 428058
rect 138954 392378 138986 392614
rect 139222 392378 139306 392614
rect 139542 392378 139574 392614
rect 138954 392294 139574 392378
rect 138954 392058 138986 392294
rect 139222 392058 139306 392294
rect 139542 392058 139574 392294
rect 138954 356614 139574 392058
rect 138954 356378 138986 356614
rect 139222 356378 139306 356614
rect 139542 356378 139574 356614
rect 138954 356294 139574 356378
rect 138954 356058 138986 356294
rect 139222 356058 139306 356294
rect 139542 356058 139574 356294
rect 138954 320614 139574 356058
rect 138954 320378 138986 320614
rect 139222 320378 139306 320614
rect 139542 320378 139574 320614
rect 138954 320294 139574 320378
rect 138954 320058 138986 320294
rect 139222 320058 139306 320294
rect 139542 320058 139574 320294
rect 138954 284614 139574 320058
rect 138954 284378 138986 284614
rect 139222 284378 139306 284614
rect 139542 284378 139574 284614
rect 138954 284294 139574 284378
rect 138954 284058 138986 284294
rect 139222 284058 139306 284294
rect 139542 284058 139574 284294
rect 138954 248614 139574 284058
rect 138954 248378 138986 248614
rect 139222 248378 139306 248614
rect 139542 248378 139574 248614
rect 138954 248294 139574 248378
rect 138954 248058 138986 248294
rect 139222 248058 139306 248294
rect 139542 248058 139574 248294
rect 138954 212614 139574 248058
rect 138954 212378 138986 212614
rect 139222 212378 139306 212614
rect 139542 212378 139574 212614
rect 138954 212294 139574 212378
rect 138954 212058 138986 212294
rect 139222 212058 139306 212294
rect 139542 212058 139574 212294
rect 138954 176614 139574 212058
rect 138954 176378 138986 176614
rect 139222 176378 139306 176614
rect 139542 176378 139574 176614
rect 138954 176294 139574 176378
rect 138954 176058 138986 176294
rect 139222 176058 139306 176294
rect 139542 176058 139574 176294
rect 138954 140614 139574 176058
rect 138954 140378 138986 140614
rect 139222 140378 139306 140614
rect 139542 140378 139574 140614
rect 138954 140294 139574 140378
rect 138954 140058 138986 140294
rect 139222 140058 139306 140294
rect 139542 140058 139574 140294
rect 138954 104614 139574 140058
rect 138954 104378 138986 104614
rect 139222 104378 139306 104614
rect 139542 104378 139574 104614
rect 138954 104294 139574 104378
rect 138954 104058 138986 104294
rect 139222 104058 139306 104294
rect 139542 104058 139574 104294
rect 138954 68614 139574 104058
rect 138954 68378 138986 68614
rect 139222 68378 139306 68614
rect 139542 68378 139574 68614
rect 138954 68294 139574 68378
rect 138954 68058 138986 68294
rect 139222 68058 139306 68294
rect 139542 68058 139574 68294
rect 138954 32614 139574 68058
rect 138954 32378 138986 32614
rect 139222 32378 139306 32614
rect 139542 32378 139574 32614
rect 138954 32294 139574 32378
rect 138954 32058 138986 32294
rect 139222 32058 139306 32294
rect 139542 32058 139574 32294
rect 120954 -6342 120986 -6106
rect 121222 -6342 121306 -6106
rect 121542 -6342 121574 -6106
rect 120954 -6426 121574 -6342
rect 120954 -6662 120986 -6426
rect 121222 -6662 121306 -6426
rect 121542 -6662 121574 -6426
rect 120954 -7654 121574 -6662
rect 138954 -7066 139574 32058
rect 145794 704838 146414 705830
rect 145794 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 146414 704838
rect 145794 704518 146414 704602
rect 145794 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 146414 704518
rect 145794 687454 146414 704282
rect 145794 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 146414 687454
rect 145794 687134 146414 687218
rect 145794 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 146414 687134
rect 145794 651454 146414 686898
rect 145794 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 146414 651454
rect 145794 651134 146414 651218
rect 145794 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 146414 651134
rect 145794 615454 146414 650898
rect 145794 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 146414 615454
rect 145794 615134 146414 615218
rect 145794 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 146414 615134
rect 145794 579454 146414 614898
rect 145794 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 146414 579454
rect 145794 579134 146414 579218
rect 145794 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 146414 579134
rect 145794 543454 146414 578898
rect 145794 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 146414 543454
rect 145794 543134 146414 543218
rect 145794 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 146414 543134
rect 145794 507454 146414 542898
rect 145794 507218 145826 507454
rect 146062 507218 146146 507454
rect 146382 507218 146414 507454
rect 145794 507134 146414 507218
rect 145794 506898 145826 507134
rect 146062 506898 146146 507134
rect 146382 506898 146414 507134
rect 145794 471454 146414 506898
rect 145794 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 146414 471454
rect 145794 471134 146414 471218
rect 145794 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 146414 471134
rect 145794 435454 146414 470898
rect 145794 435218 145826 435454
rect 146062 435218 146146 435454
rect 146382 435218 146414 435454
rect 145794 435134 146414 435218
rect 145794 434898 145826 435134
rect 146062 434898 146146 435134
rect 146382 434898 146414 435134
rect 145794 399454 146414 434898
rect 145794 399218 145826 399454
rect 146062 399218 146146 399454
rect 146382 399218 146414 399454
rect 145794 399134 146414 399218
rect 145794 398898 145826 399134
rect 146062 398898 146146 399134
rect 146382 398898 146414 399134
rect 145794 363454 146414 398898
rect 145794 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 146414 363454
rect 145794 363134 146414 363218
rect 145794 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 146414 363134
rect 145794 327454 146414 362898
rect 145794 327218 145826 327454
rect 146062 327218 146146 327454
rect 146382 327218 146414 327454
rect 145794 327134 146414 327218
rect 145794 326898 145826 327134
rect 146062 326898 146146 327134
rect 146382 326898 146414 327134
rect 145794 291454 146414 326898
rect 145794 291218 145826 291454
rect 146062 291218 146146 291454
rect 146382 291218 146414 291454
rect 145794 291134 146414 291218
rect 145794 290898 145826 291134
rect 146062 290898 146146 291134
rect 146382 290898 146414 291134
rect 145794 255454 146414 290898
rect 145794 255218 145826 255454
rect 146062 255218 146146 255454
rect 146382 255218 146414 255454
rect 145794 255134 146414 255218
rect 145794 254898 145826 255134
rect 146062 254898 146146 255134
rect 146382 254898 146414 255134
rect 145794 219454 146414 254898
rect 145794 219218 145826 219454
rect 146062 219218 146146 219454
rect 146382 219218 146414 219454
rect 145794 219134 146414 219218
rect 145794 218898 145826 219134
rect 146062 218898 146146 219134
rect 146382 218898 146414 219134
rect 145794 183454 146414 218898
rect 145794 183218 145826 183454
rect 146062 183218 146146 183454
rect 146382 183218 146414 183454
rect 145794 183134 146414 183218
rect 145794 182898 145826 183134
rect 146062 182898 146146 183134
rect 146382 182898 146414 183134
rect 145794 147454 146414 182898
rect 145794 147218 145826 147454
rect 146062 147218 146146 147454
rect 146382 147218 146414 147454
rect 145794 147134 146414 147218
rect 145794 146898 145826 147134
rect 146062 146898 146146 147134
rect 146382 146898 146414 147134
rect 145794 111454 146414 146898
rect 145794 111218 145826 111454
rect 146062 111218 146146 111454
rect 146382 111218 146414 111454
rect 145794 111134 146414 111218
rect 145794 110898 145826 111134
rect 146062 110898 146146 111134
rect 146382 110898 146414 111134
rect 145794 75454 146414 110898
rect 145794 75218 145826 75454
rect 146062 75218 146146 75454
rect 146382 75218 146414 75454
rect 145794 75134 146414 75218
rect 145794 74898 145826 75134
rect 146062 74898 146146 75134
rect 146382 74898 146414 75134
rect 145794 39454 146414 74898
rect 145794 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 146414 39454
rect 145794 39134 146414 39218
rect 145794 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 146414 39134
rect 145794 3454 146414 38898
rect 145794 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 146414 3454
rect 145794 3134 146414 3218
rect 145794 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 146414 3134
rect 145794 -346 146414 2898
rect 145794 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 146414 -346
rect 145794 -666 146414 -582
rect 145794 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 146414 -666
rect 145794 -1894 146414 -902
rect 149514 691174 150134 706202
rect 149514 690938 149546 691174
rect 149782 690938 149866 691174
rect 150102 690938 150134 691174
rect 149514 690854 150134 690938
rect 149514 690618 149546 690854
rect 149782 690618 149866 690854
rect 150102 690618 150134 690854
rect 149514 655174 150134 690618
rect 149514 654938 149546 655174
rect 149782 654938 149866 655174
rect 150102 654938 150134 655174
rect 149514 654854 150134 654938
rect 149514 654618 149546 654854
rect 149782 654618 149866 654854
rect 150102 654618 150134 654854
rect 149514 619174 150134 654618
rect 149514 618938 149546 619174
rect 149782 618938 149866 619174
rect 150102 618938 150134 619174
rect 149514 618854 150134 618938
rect 149514 618618 149546 618854
rect 149782 618618 149866 618854
rect 150102 618618 150134 618854
rect 149514 583174 150134 618618
rect 149514 582938 149546 583174
rect 149782 582938 149866 583174
rect 150102 582938 150134 583174
rect 149514 582854 150134 582938
rect 149514 582618 149546 582854
rect 149782 582618 149866 582854
rect 150102 582618 150134 582854
rect 149514 547174 150134 582618
rect 149514 546938 149546 547174
rect 149782 546938 149866 547174
rect 150102 546938 150134 547174
rect 149514 546854 150134 546938
rect 149514 546618 149546 546854
rect 149782 546618 149866 546854
rect 150102 546618 150134 546854
rect 149514 511174 150134 546618
rect 149514 510938 149546 511174
rect 149782 510938 149866 511174
rect 150102 510938 150134 511174
rect 149514 510854 150134 510938
rect 149514 510618 149546 510854
rect 149782 510618 149866 510854
rect 150102 510618 150134 510854
rect 149514 475174 150134 510618
rect 149514 474938 149546 475174
rect 149782 474938 149866 475174
rect 150102 474938 150134 475174
rect 149514 474854 150134 474938
rect 149514 474618 149546 474854
rect 149782 474618 149866 474854
rect 150102 474618 150134 474854
rect 149514 439174 150134 474618
rect 149514 438938 149546 439174
rect 149782 438938 149866 439174
rect 150102 438938 150134 439174
rect 149514 438854 150134 438938
rect 149514 438618 149546 438854
rect 149782 438618 149866 438854
rect 150102 438618 150134 438854
rect 149514 403174 150134 438618
rect 149514 402938 149546 403174
rect 149782 402938 149866 403174
rect 150102 402938 150134 403174
rect 149514 402854 150134 402938
rect 149514 402618 149546 402854
rect 149782 402618 149866 402854
rect 150102 402618 150134 402854
rect 149514 367174 150134 402618
rect 149514 366938 149546 367174
rect 149782 366938 149866 367174
rect 150102 366938 150134 367174
rect 149514 366854 150134 366938
rect 149514 366618 149546 366854
rect 149782 366618 149866 366854
rect 150102 366618 150134 366854
rect 149514 331174 150134 366618
rect 149514 330938 149546 331174
rect 149782 330938 149866 331174
rect 150102 330938 150134 331174
rect 149514 330854 150134 330938
rect 149514 330618 149546 330854
rect 149782 330618 149866 330854
rect 150102 330618 150134 330854
rect 149514 295174 150134 330618
rect 149514 294938 149546 295174
rect 149782 294938 149866 295174
rect 150102 294938 150134 295174
rect 149514 294854 150134 294938
rect 149514 294618 149546 294854
rect 149782 294618 149866 294854
rect 150102 294618 150134 294854
rect 149514 259174 150134 294618
rect 149514 258938 149546 259174
rect 149782 258938 149866 259174
rect 150102 258938 150134 259174
rect 149514 258854 150134 258938
rect 149514 258618 149546 258854
rect 149782 258618 149866 258854
rect 150102 258618 150134 258854
rect 149514 223174 150134 258618
rect 149514 222938 149546 223174
rect 149782 222938 149866 223174
rect 150102 222938 150134 223174
rect 149514 222854 150134 222938
rect 149514 222618 149546 222854
rect 149782 222618 149866 222854
rect 150102 222618 150134 222854
rect 149514 187174 150134 222618
rect 149514 186938 149546 187174
rect 149782 186938 149866 187174
rect 150102 186938 150134 187174
rect 149514 186854 150134 186938
rect 149514 186618 149546 186854
rect 149782 186618 149866 186854
rect 150102 186618 150134 186854
rect 149514 151174 150134 186618
rect 149514 150938 149546 151174
rect 149782 150938 149866 151174
rect 150102 150938 150134 151174
rect 149514 150854 150134 150938
rect 149514 150618 149546 150854
rect 149782 150618 149866 150854
rect 150102 150618 150134 150854
rect 149514 115174 150134 150618
rect 149514 114938 149546 115174
rect 149782 114938 149866 115174
rect 150102 114938 150134 115174
rect 149514 114854 150134 114938
rect 149514 114618 149546 114854
rect 149782 114618 149866 114854
rect 150102 114618 150134 114854
rect 149514 79174 150134 114618
rect 149514 78938 149546 79174
rect 149782 78938 149866 79174
rect 150102 78938 150134 79174
rect 149514 78854 150134 78938
rect 149514 78618 149546 78854
rect 149782 78618 149866 78854
rect 150102 78618 150134 78854
rect 149514 43174 150134 78618
rect 149514 42938 149546 43174
rect 149782 42938 149866 43174
rect 150102 42938 150134 43174
rect 149514 42854 150134 42938
rect 149514 42618 149546 42854
rect 149782 42618 149866 42854
rect 150102 42618 150134 42854
rect 149514 7174 150134 42618
rect 149514 6938 149546 7174
rect 149782 6938 149866 7174
rect 150102 6938 150134 7174
rect 149514 6854 150134 6938
rect 149514 6618 149546 6854
rect 149782 6618 149866 6854
rect 150102 6618 150134 6854
rect 149514 -2266 150134 6618
rect 149514 -2502 149546 -2266
rect 149782 -2502 149866 -2266
rect 150102 -2502 150134 -2266
rect 149514 -2586 150134 -2502
rect 149514 -2822 149546 -2586
rect 149782 -2822 149866 -2586
rect 150102 -2822 150134 -2586
rect 149514 -3814 150134 -2822
rect 153234 694894 153854 708122
rect 153234 694658 153266 694894
rect 153502 694658 153586 694894
rect 153822 694658 153854 694894
rect 153234 694574 153854 694658
rect 153234 694338 153266 694574
rect 153502 694338 153586 694574
rect 153822 694338 153854 694574
rect 153234 658894 153854 694338
rect 153234 658658 153266 658894
rect 153502 658658 153586 658894
rect 153822 658658 153854 658894
rect 153234 658574 153854 658658
rect 153234 658338 153266 658574
rect 153502 658338 153586 658574
rect 153822 658338 153854 658574
rect 153234 622894 153854 658338
rect 153234 622658 153266 622894
rect 153502 622658 153586 622894
rect 153822 622658 153854 622894
rect 153234 622574 153854 622658
rect 153234 622338 153266 622574
rect 153502 622338 153586 622574
rect 153822 622338 153854 622574
rect 153234 586894 153854 622338
rect 153234 586658 153266 586894
rect 153502 586658 153586 586894
rect 153822 586658 153854 586894
rect 153234 586574 153854 586658
rect 153234 586338 153266 586574
rect 153502 586338 153586 586574
rect 153822 586338 153854 586574
rect 153234 550894 153854 586338
rect 153234 550658 153266 550894
rect 153502 550658 153586 550894
rect 153822 550658 153854 550894
rect 153234 550574 153854 550658
rect 153234 550338 153266 550574
rect 153502 550338 153586 550574
rect 153822 550338 153854 550574
rect 153234 514894 153854 550338
rect 153234 514658 153266 514894
rect 153502 514658 153586 514894
rect 153822 514658 153854 514894
rect 153234 514574 153854 514658
rect 153234 514338 153266 514574
rect 153502 514338 153586 514574
rect 153822 514338 153854 514574
rect 153234 478894 153854 514338
rect 153234 478658 153266 478894
rect 153502 478658 153586 478894
rect 153822 478658 153854 478894
rect 153234 478574 153854 478658
rect 153234 478338 153266 478574
rect 153502 478338 153586 478574
rect 153822 478338 153854 478574
rect 153234 442894 153854 478338
rect 153234 442658 153266 442894
rect 153502 442658 153586 442894
rect 153822 442658 153854 442894
rect 153234 442574 153854 442658
rect 153234 442338 153266 442574
rect 153502 442338 153586 442574
rect 153822 442338 153854 442574
rect 153234 406894 153854 442338
rect 153234 406658 153266 406894
rect 153502 406658 153586 406894
rect 153822 406658 153854 406894
rect 153234 406574 153854 406658
rect 153234 406338 153266 406574
rect 153502 406338 153586 406574
rect 153822 406338 153854 406574
rect 153234 370894 153854 406338
rect 153234 370658 153266 370894
rect 153502 370658 153586 370894
rect 153822 370658 153854 370894
rect 153234 370574 153854 370658
rect 153234 370338 153266 370574
rect 153502 370338 153586 370574
rect 153822 370338 153854 370574
rect 153234 334894 153854 370338
rect 153234 334658 153266 334894
rect 153502 334658 153586 334894
rect 153822 334658 153854 334894
rect 153234 334574 153854 334658
rect 153234 334338 153266 334574
rect 153502 334338 153586 334574
rect 153822 334338 153854 334574
rect 153234 298894 153854 334338
rect 153234 298658 153266 298894
rect 153502 298658 153586 298894
rect 153822 298658 153854 298894
rect 153234 298574 153854 298658
rect 153234 298338 153266 298574
rect 153502 298338 153586 298574
rect 153822 298338 153854 298574
rect 153234 262894 153854 298338
rect 153234 262658 153266 262894
rect 153502 262658 153586 262894
rect 153822 262658 153854 262894
rect 153234 262574 153854 262658
rect 153234 262338 153266 262574
rect 153502 262338 153586 262574
rect 153822 262338 153854 262574
rect 153234 226894 153854 262338
rect 153234 226658 153266 226894
rect 153502 226658 153586 226894
rect 153822 226658 153854 226894
rect 153234 226574 153854 226658
rect 153234 226338 153266 226574
rect 153502 226338 153586 226574
rect 153822 226338 153854 226574
rect 153234 190894 153854 226338
rect 153234 190658 153266 190894
rect 153502 190658 153586 190894
rect 153822 190658 153854 190894
rect 153234 190574 153854 190658
rect 153234 190338 153266 190574
rect 153502 190338 153586 190574
rect 153822 190338 153854 190574
rect 153234 154894 153854 190338
rect 153234 154658 153266 154894
rect 153502 154658 153586 154894
rect 153822 154658 153854 154894
rect 153234 154574 153854 154658
rect 153234 154338 153266 154574
rect 153502 154338 153586 154574
rect 153822 154338 153854 154574
rect 153234 118894 153854 154338
rect 153234 118658 153266 118894
rect 153502 118658 153586 118894
rect 153822 118658 153854 118894
rect 153234 118574 153854 118658
rect 153234 118338 153266 118574
rect 153502 118338 153586 118574
rect 153822 118338 153854 118574
rect 153234 82894 153854 118338
rect 153234 82658 153266 82894
rect 153502 82658 153586 82894
rect 153822 82658 153854 82894
rect 153234 82574 153854 82658
rect 153234 82338 153266 82574
rect 153502 82338 153586 82574
rect 153822 82338 153854 82574
rect 153234 46894 153854 82338
rect 153234 46658 153266 46894
rect 153502 46658 153586 46894
rect 153822 46658 153854 46894
rect 153234 46574 153854 46658
rect 153234 46338 153266 46574
rect 153502 46338 153586 46574
rect 153822 46338 153854 46574
rect 153234 10894 153854 46338
rect 153234 10658 153266 10894
rect 153502 10658 153586 10894
rect 153822 10658 153854 10894
rect 153234 10574 153854 10658
rect 153234 10338 153266 10574
rect 153502 10338 153586 10574
rect 153822 10338 153854 10574
rect 153234 -4186 153854 10338
rect 153234 -4422 153266 -4186
rect 153502 -4422 153586 -4186
rect 153822 -4422 153854 -4186
rect 153234 -4506 153854 -4422
rect 153234 -4742 153266 -4506
rect 153502 -4742 153586 -4506
rect 153822 -4742 153854 -4506
rect 153234 -5734 153854 -4742
rect 156954 698614 157574 710042
rect 174954 711558 175574 711590
rect 174954 711322 174986 711558
rect 175222 711322 175306 711558
rect 175542 711322 175574 711558
rect 174954 711238 175574 711322
rect 174954 711002 174986 711238
rect 175222 711002 175306 711238
rect 175542 711002 175574 711238
rect 171234 709638 171854 709670
rect 171234 709402 171266 709638
rect 171502 709402 171586 709638
rect 171822 709402 171854 709638
rect 171234 709318 171854 709402
rect 171234 709082 171266 709318
rect 171502 709082 171586 709318
rect 171822 709082 171854 709318
rect 167514 707718 168134 707750
rect 167514 707482 167546 707718
rect 167782 707482 167866 707718
rect 168102 707482 168134 707718
rect 167514 707398 168134 707482
rect 167514 707162 167546 707398
rect 167782 707162 167866 707398
rect 168102 707162 168134 707398
rect 156954 698378 156986 698614
rect 157222 698378 157306 698614
rect 157542 698378 157574 698614
rect 156954 698294 157574 698378
rect 156954 698058 156986 698294
rect 157222 698058 157306 698294
rect 157542 698058 157574 698294
rect 156954 662614 157574 698058
rect 156954 662378 156986 662614
rect 157222 662378 157306 662614
rect 157542 662378 157574 662614
rect 156954 662294 157574 662378
rect 156954 662058 156986 662294
rect 157222 662058 157306 662294
rect 157542 662058 157574 662294
rect 156954 626614 157574 662058
rect 156954 626378 156986 626614
rect 157222 626378 157306 626614
rect 157542 626378 157574 626614
rect 156954 626294 157574 626378
rect 156954 626058 156986 626294
rect 157222 626058 157306 626294
rect 157542 626058 157574 626294
rect 156954 590614 157574 626058
rect 156954 590378 156986 590614
rect 157222 590378 157306 590614
rect 157542 590378 157574 590614
rect 156954 590294 157574 590378
rect 156954 590058 156986 590294
rect 157222 590058 157306 590294
rect 157542 590058 157574 590294
rect 156954 554614 157574 590058
rect 156954 554378 156986 554614
rect 157222 554378 157306 554614
rect 157542 554378 157574 554614
rect 156954 554294 157574 554378
rect 156954 554058 156986 554294
rect 157222 554058 157306 554294
rect 157542 554058 157574 554294
rect 156954 518614 157574 554058
rect 156954 518378 156986 518614
rect 157222 518378 157306 518614
rect 157542 518378 157574 518614
rect 156954 518294 157574 518378
rect 156954 518058 156986 518294
rect 157222 518058 157306 518294
rect 157542 518058 157574 518294
rect 156954 482614 157574 518058
rect 163794 705798 164414 705830
rect 163794 705562 163826 705798
rect 164062 705562 164146 705798
rect 164382 705562 164414 705798
rect 163794 705478 164414 705562
rect 163794 705242 163826 705478
rect 164062 705242 164146 705478
rect 164382 705242 164414 705478
rect 163794 669454 164414 705242
rect 163794 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 164414 669454
rect 163794 669134 164414 669218
rect 163794 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 164414 669134
rect 163794 633454 164414 668898
rect 163794 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 164414 633454
rect 163794 633134 164414 633218
rect 163794 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 164414 633134
rect 163794 597454 164414 632898
rect 163794 597218 163826 597454
rect 164062 597218 164146 597454
rect 164382 597218 164414 597454
rect 163794 597134 164414 597218
rect 163794 596898 163826 597134
rect 164062 596898 164146 597134
rect 164382 596898 164414 597134
rect 163794 561454 164414 596898
rect 163794 561218 163826 561454
rect 164062 561218 164146 561454
rect 164382 561218 164414 561454
rect 163794 561134 164414 561218
rect 163794 560898 163826 561134
rect 164062 560898 164146 561134
rect 164382 560898 164414 561134
rect 163794 525454 164414 560898
rect 163794 525218 163826 525454
rect 164062 525218 164146 525454
rect 164382 525218 164414 525454
rect 163794 525134 164414 525218
rect 163794 524898 163826 525134
rect 164062 524898 164146 525134
rect 164382 524898 164414 525134
rect 163794 509939 164414 524898
rect 167514 673174 168134 707162
rect 167514 672938 167546 673174
rect 167782 672938 167866 673174
rect 168102 672938 168134 673174
rect 167514 672854 168134 672938
rect 167514 672618 167546 672854
rect 167782 672618 167866 672854
rect 168102 672618 168134 672854
rect 167514 637174 168134 672618
rect 167514 636938 167546 637174
rect 167782 636938 167866 637174
rect 168102 636938 168134 637174
rect 167514 636854 168134 636938
rect 167514 636618 167546 636854
rect 167782 636618 167866 636854
rect 168102 636618 168134 636854
rect 167514 601174 168134 636618
rect 167514 600938 167546 601174
rect 167782 600938 167866 601174
rect 168102 600938 168134 601174
rect 167514 600854 168134 600938
rect 167514 600618 167546 600854
rect 167782 600618 167866 600854
rect 168102 600618 168134 600854
rect 167514 565174 168134 600618
rect 167514 564938 167546 565174
rect 167782 564938 167866 565174
rect 168102 564938 168134 565174
rect 167514 564854 168134 564938
rect 167514 564618 167546 564854
rect 167782 564618 167866 564854
rect 168102 564618 168134 564854
rect 167514 529174 168134 564618
rect 167514 528938 167546 529174
rect 167782 528938 167866 529174
rect 168102 528938 168134 529174
rect 167514 528854 168134 528938
rect 167514 528618 167546 528854
rect 167782 528618 167866 528854
rect 168102 528618 168134 528854
rect 167514 509939 168134 528618
rect 171234 676894 171854 709082
rect 171234 676658 171266 676894
rect 171502 676658 171586 676894
rect 171822 676658 171854 676894
rect 171234 676574 171854 676658
rect 171234 676338 171266 676574
rect 171502 676338 171586 676574
rect 171822 676338 171854 676574
rect 171234 640894 171854 676338
rect 171234 640658 171266 640894
rect 171502 640658 171586 640894
rect 171822 640658 171854 640894
rect 171234 640574 171854 640658
rect 171234 640338 171266 640574
rect 171502 640338 171586 640574
rect 171822 640338 171854 640574
rect 171234 604894 171854 640338
rect 171234 604658 171266 604894
rect 171502 604658 171586 604894
rect 171822 604658 171854 604894
rect 171234 604574 171854 604658
rect 171234 604338 171266 604574
rect 171502 604338 171586 604574
rect 171822 604338 171854 604574
rect 171234 568894 171854 604338
rect 171234 568658 171266 568894
rect 171502 568658 171586 568894
rect 171822 568658 171854 568894
rect 171234 568574 171854 568658
rect 171234 568338 171266 568574
rect 171502 568338 171586 568574
rect 171822 568338 171854 568574
rect 171234 532894 171854 568338
rect 171234 532658 171266 532894
rect 171502 532658 171586 532894
rect 171822 532658 171854 532894
rect 171234 532574 171854 532658
rect 171234 532338 171266 532574
rect 171502 532338 171586 532574
rect 171822 532338 171854 532574
rect 171234 509939 171854 532338
rect 174954 680614 175574 711002
rect 192954 710598 193574 711590
rect 192954 710362 192986 710598
rect 193222 710362 193306 710598
rect 193542 710362 193574 710598
rect 192954 710278 193574 710362
rect 192954 710042 192986 710278
rect 193222 710042 193306 710278
rect 193542 710042 193574 710278
rect 189234 708678 189854 709670
rect 189234 708442 189266 708678
rect 189502 708442 189586 708678
rect 189822 708442 189854 708678
rect 189234 708358 189854 708442
rect 189234 708122 189266 708358
rect 189502 708122 189586 708358
rect 189822 708122 189854 708358
rect 185514 706758 186134 707750
rect 185514 706522 185546 706758
rect 185782 706522 185866 706758
rect 186102 706522 186134 706758
rect 185514 706438 186134 706522
rect 185514 706202 185546 706438
rect 185782 706202 185866 706438
rect 186102 706202 186134 706438
rect 174954 680378 174986 680614
rect 175222 680378 175306 680614
rect 175542 680378 175574 680614
rect 174954 680294 175574 680378
rect 174954 680058 174986 680294
rect 175222 680058 175306 680294
rect 175542 680058 175574 680294
rect 174954 644614 175574 680058
rect 174954 644378 174986 644614
rect 175222 644378 175306 644614
rect 175542 644378 175574 644614
rect 174954 644294 175574 644378
rect 174954 644058 174986 644294
rect 175222 644058 175306 644294
rect 175542 644058 175574 644294
rect 174954 608614 175574 644058
rect 174954 608378 174986 608614
rect 175222 608378 175306 608614
rect 175542 608378 175574 608614
rect 174954 608294 175574 608378
rect 174954 608058 174986 608294
rect 175222 608058 175306 608294
rect 175542 608058 175574 608294
rect 174954 572614 175574 608058
rect 174954 572378 174986 572614
rect 175222 572378 175306 572614
rect 175542 572378 175574 572614
rect 174954 572294 175574 572378
rect 174954 572058 174986 572294
rect 175222 572058 175306 572294
rect 175542 572058 175574 572294
rect 174954 536614 175574 572058
rect 174954 536378 174986 536614
rect 175222 536378 175306 536614
rect 175542 536378 175574 536614
rect 174954 536294 175574 536378
rect 174954 536058 174986 536294
rect 175222 536058 175306 536294
rect 175542 536058 175574 536294
rect 174954 509939 175574 536058
rect 181794 704838 182414 705830
rect 181794 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 182414 704838
rect 181794 704518 182414 704602
rect 181794 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 182414 704518
rect 181794 687454 182414 704282
rect 181794 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 182414 687454
rect 181794 687134 182414 687218
rect 181794 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 182414 687134
rect 181794 651454 182414 686898
rect 181794 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 182414 651454
rect 181794 651134 182414 651218
rect 181794 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 182414 651134
rect 181794 615454 182414 650898
rect 181794 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 182414 615454
rect 181794 615134 182414 615218
rect 181794 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 182414 615134
rect 181794 579454 182414 614898
rect 181794 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 182414 579454
rect 181794 579134 182414 579218
rect 181794 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 182414 579134
rect 181794 543454 182414 578898
rect 181794 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 182414 543454
rect 181794 543134 182414 543218
rect 181794 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 182414 543134
rect 181794 509939 182414 542898
rect 185514 691174 186134 706202
rect 185514 690938 185546 691174
rect 185782 690938 185866 691174
rect 186102 690938 186134 691174
rect 185514 690854 186134 690938
rect 185514 690618 185546 690854
rect 185782 690618 185866 690854
rect 186102 690618 186134 690854
rect 185514 655174 186134 690618
rect 185514 654938 185546 655174
rect 185782 654938 185866 655174
rect 186102 654938 186134 655174
rect 185514 654854 186134 654938
rect 185514 654618 185546 654854
rect 185782 654618 185866 654854
rect 186102 654618 186134 654854
rect 185514 619174 186134 654618
rect 185514 618938 185546 619174
rect 185782 618938 185866 619174
rect 186102 618938 186134 619174
rect 185514 618854 186134 618938
rect 185514 618618 185546 618854
rect 185782 618618 185866 618854
rect 186102 618618 186134 618854
rect 185514 583174 186134 618618
rect 185514 582938 185546 583174
rect 185782 582938 185866 583174
rect 186102 582938 186134 583174
rect 185514 582854 186134 582938
rect 185514 582618 185546 582854
rect 185782 582618 185866 582854
rect 186102 582618 186134 582854
rect 185514 547174 186134 582618
rect 185514 546938 185546 547174
rect 185782 546938 185866 547174
rect 186102 546938 186134 547174
rect 185514 546854 186134 546938
rect 185514 546618 185546 546854
rect 185782 546618 185866 546854
rect 186102 546618 186134 546854
rect 185514 511174 186134 546618
rect 185514 510938 185546 511174
rect 185782 510938 185866 511174
rect 186102 510938 186134 511174
rect 185514 510854 186134 510938
rect 185514 510618 185546 510854
rect 185782 510618 185866 510854
rect 186102 510618 186134 510854
rect 185514 509939 186134 510618
rect 189234 694894 189854 708122
rect 189234 694658 189266 694894
rect 189502 694658 189586 694894
rect 189822 694658 189854 694894
rect 189234 694574 189854 694658
rect 189234 694338 189266 694574
rect 189502 694338 189586 694574
rect 189822 694338 189854 694574
rect 189234 658894 189854 694338
rect 189234 658658 189266 658894
rect 189502 658658 189586 658894
rect 189822 658658 189854 658894
rect 189234 658574 189854 658658
rect 189234 658338 189266 658574
rect 189502 658338 189586 658574
rect 189822 658338 189854 658574
rect 189234 622894 189854 658338
rect 189234 622658 189266 622894
rect 189502 622658 189586 622894
rect 189822 622658 189854 622894
rect 189234 622574 189854 622658
rect 189234 622338 189266 622574
rect 189502 622338 189586 622574
rect 189822 622338 189854 622574
rect 189234 586894 189854 622338
rect 189234 586658 189266 586894
rect 189502 586658 189586 586894
rect 189822 586658 189854 586894
rect 189234 586574 189854 586658
rect 189234 586338 189266 586574
rect 189502 586338 189586 586574
rect 189822 586338 189854 586574
rect 189234 550894 189854 586338
rect 189234 550658 189266 550894
rect 189502 550658 189586 550894
rect 189822 550658 189854 550894
rect 189234 550574 189854 550658
rect 189234 550338 189266 550574
rect 189502 550338 189586 550574
rect 189822 550338 189854 550574
rect 189234 514894 189854 550338
rect 189234 514658 189266 514894
rect 189502 514658 189586 514894
rect 189822 514658 189854 514894
rect 189234 514574 189854 514658
rect 189234 514338 189266 514574
rect 189502 514338 189586 514574
rect 189822 514338 189854 514574
rect 189234 509939 189854 514338
rect 192954 698614 193574 710042
rect 210954 711558 211574 711590
rect 210954 711322 210986 711558
rect 211222 711322 211306 711558
rect 211542 711322 211574 711558
rect 210954 711238 211574 711322
rect 210954 711002 210986 711238
rect 211222 711002 211306 711238
rect 211542 711002 211574 711238
rect 207234 709638 207854 709670
rect 207234 709402 207266 709638
rect 207502 709402 207586 709638
rect 207822 709402 207854 709638
rect 207234 709318 207854 709402
rect 207234 709082 207266 709318
rect 207502 709082 207586 709318
rect 207822 709082 207854 709318
rect 203514 707718 204134 707750
rect 203514 707482 203546 707718
rect 203782 707482 203866 707718
rect 204102 707482 204134 707718
rect 203514 707398 204134 707482
rect 203514 707162 203546 707398
rect 203782 707162 203866 707398
rect 204102 707162 204134 707398
rect 192954 698378 192986 698614
rect 193222 698378 193306 698614
rect 193542 698378 193574 698614
rect 192954 698294 193574 698378
rect 192954 698058 192986 698294
rect 193222 698058 193306 698294
rect 193542 698058 193574 698294
rect 192954 662614 193574 698058
rect 192954 662378 192986 662614
rect 193222 662378 193306 662614
rect 193542 662378 193574 662614
rect 192954 662294 193574 662378
rect 192954 662058 192986 662294
rect 193222 662058 193306 662294
rect 193542 662058 193574 662294
rect 192954 626614 193574 662058
rect 192954 626378 192986 626614
rect 193222 626378 193306 626614
rect 193542 626378 193574 626614
rect 192954 626294 193574 626378
rect 192954 626058 192986 626294
rect 193222 626058 193306 626294
rect 193542 626058 193574 626294
rect 192954 590614 193574 626058
rect 192954 590378 192986 590614
rect 193222 590378 193306 590614
rect 193542 590378 193574 590614
rect 192954 590294 193574 590378
rect 192954 590058 192986 590294
rect 193222 590058 193306 590294
rect 193542 590058 193574 590294
rect 192954 554614 193574 590058
rect 192954 554378 192986 554614
rect 193222 554378 193306 554614
rect 193542 554378 193574 554614
rect 192954 554294 193574 554378
rect 192954 554058 192986 554294
rect 193222 554058 193306 554294
rect 193542 554058 193574 554294
rect 192954 518614 193574 554058
rect 192954 518378 192986 518614
rect 193222 518378 193306 518614
rect 193542 518378 193574 518614
rect 192954 518294 193574 518378
rect 192954 518058 192986 518294
rect 193222 518058 193306 518294
rect 193542 518058 193574 518294
rect 192954 509939 193574 518058
rect 199794 705798 200414 705830
rect 199794 705562 199826 705798
rect 200062 705562 200146 705798
rect 200382 705562 200414 705798
rect 199794 705478 200414 705562
rect 199794 705242 199826 705478
rect 200062 705242 200146 705478
rect 200382 705242 200414 705478
rect 199794 669454 200414 705242
rect 199794 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 200414 669454
rect 199794 669134 200414 669218
rect 199794 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 200414 669134
rect 199794 633454 200414 668898
rect 199794 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 200414 633454
rect 199794 633134 200414 633218
rect 199794 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 200414 633134
rect 199794 597454 200414 632898
rect 199794 597218 199826 597454
rect 200062 597218 200146 597454
rect 200382 597218 200414 597454
rect 199794 597134 200414 597218
rect 199794 596898 199826 597134
rect 200062 596898 200146 597134
rect 200382 596898 200414 597134
rect 199794 561454 200414 596898
rect 199794 561218 199826 561454
rect 200062 561218 200146 561454
rect 200382 561218 200414 561454
rect 199794 561134 200414 561218
rect 199794 560898 199826 561134
rect 200062 560898 200146 561134
rect 200382 560898 200414 561134
rect 199794 525454 200414 560898
rect 199794 525218 199826 525454
rect 200062 525218 200146 525454
rect 200382 525218 200414 525454
rect 199794 525134 200414 525218
rect 199794 524898 199826 525134
rect 200062 524898 200146 525134
rect 200382 524898 200414 525134
rect 199794 509939 200414 524898
rect 203514 673174 204134 707162
rect 203514 672938 203546 673174
rect 203782 672938 203866 673174
rect 204102 672938 204134 673174
rect 203514 672854 204134 672938
rect 203514 672618 203546 672854
rect 203782 672618 203866 672854
rect 204102 672618 204134 672854
rect 203514 637174 204134 672618
rect 203514 636938 203546 637174
rect 203782 636938 203866 637174
rect 204102 636938 204134 637174
rect 203514 636854 204134 636938
rect 203514 636618 203546 636854
rect 203782 636618 203866 636854
rect 204102 636618 204134 636854
rect 203514 601174 204134 636618
rect 203514 600938 203546 601174
rect 203782 600938 203866 601174
rect 204102 600938 204134 601174
rect 203514 600854 204134 600938
rect 203514 600618 203546 600854
rect 203782 600618 203866 600854
rect 204102 600618 204134 600854
rect 203514 565174 204134 600618
rect 203514 564938 203546 565174
rect 203782 564938 203866 565174
rect 204102 564938 204134 565174
rect 203514 564854 204134 564938
rect 203514 564618 203546 564854
rect 203782 564618 203866 564854
rect 204102 564618 204134 564854
rect 203514 529174 204134 564618
rect 203514 528938 203546 529174
rect 203782 528938 203866 529174
rect 204102 528938 204134 529174
rect 203514 528854 204134 528938
rect 203514 528618 203546 528854
rect 203782 528618 203866 528854
rect 204102 528618 204134 528854
rect 203514 509939 204134 528618
rect 207234 676894 207854 709082
rect 207234 676658 207266 676894
rect 207502 676658 207586 676894
rect 207822 676658 207854 676894
rect 207234 676574 207854 676658
rect 207234 676338 207266 676574
rect 207502 676338 207586 676574
rect 207822 676338 207854 676574
rect 207234 640894 207854 676338
rect 207234 640658 207266 640894
rect 207502 640658 207586 640894
rect 207822 640658 207854 640894
rect 207234 640574 207854 640658
rect 207234 640338 207266 640574
rect 207502 640338 207586 640574
rect 207822 640338 207854 640574
rect 207234 604894 207854 640338
rect 207234 604658 207266 604894
rect 207502 604658 207586 604894
rect 207822 604658 207854 604894
rect 207234 604574 207854 604658
rect 207234 604338 207266 604574
rect 207502 604338 207586 604574
rect 207822 604338 207854 604574
rect 207234 568894 207854 604338
rect 207234 568658 207266 568894
rect 207502 568658 207586 568894
rect 207822 568658 207854 568894
rect 207234 568574 207854 568658
rect 207234 568338 207266 568574
rect 207502 568338 207586 568574
rect 207822 568338 207854 568574
rect 207234 532894 207854 568338
rect 207234 532658 207266 532894
rect 207502 532658 207586 532894
rect 207822 532658 207854 532894
rect 207234 532574 207854 532658
rect 207234 532338 207266 532574
rect 207502 532338 207586 532574
rect 207822 532338 207854 532574
rect 207234 509939 207854 532338
rect 210954 680614 211574 711002
rect 228954 710598 229574 711590
rect 228954 710362 228986 710598
rect 229222 710362 229306 710598
rect 229542 710362 229574 710598
rect 228954 710278 229574 710362
rect 228954 710042 228986 710278
rect 229222 710042 229306 710278
rect 229542 710042 229574 710278
rect 225234 708678 225854 709670
rect 225234 708442 225266 708678
rect 225502 708442 225586 708678
rect 225822 708442 225854 708678
rect 225234 708358 225854 708442
rect 225234 708122 225266 708358
rect 225502 708122 225586 708358
rect 225822 708122 225854 708358
rect 221514 706758 222134 707750
rect 221514 706522 221546 706758
rect 221782 706522 221866 706758
rect 222102 706522 222134 706758
rect 221514 706438 222134 706522
rect 221514 706202 221546 706438
rect 221782 706202 221866 706438
rect 222102 706202 222134 706438
rect 210954 680378 210986 680614
rect 211222 680378 211306 680614
rect 211542 680378 211574 680614
rect 210954 680294 211574 680378
rect 210954 680058 210986 680294
rect 211222 680058 211306 680294
rect 211542 680058 211574 680294
rect 210954 644614 211574 680058
rect 210954 644378 210986 644614
rect 211222 644378 211306 644614
rect 211542 644378 211574 644614
rect 210954 644294 211574 644378
rect 210954 644058 210986 644294
rect 211222 644058 211306 644294
rect 211542 644058 211574 644294
rect 210954 608614 211574 644058
rect 210954 608378 210986 608614
rect 211222 608378 211306 608614
rect 211542 608378 211574 608614
rect 210954 608294 211574 608378
rect 210954 608058 210986 608294
rect 211222 608058 211306 608294
rect 211542 608058 211574 608294
rect 210954 572614 211574 608058
rect 210954 572378 210986 572614
rect 211222 572378 211306 572614
rect 211542 572378 211574 572614
rect 210954 572294 211574 572378
rect 210954 572058 210986 572294
rect 211222 572058 211306 572294
rect 211542 572058 211574 572294
rect 210954 536614 211574 572058
rect 210954 536378 210986 536614
rect 211222 536378 211306 536614
rect 211542 536378 211574 536614
rect 210954 536294 211574 536378
rect 210954 536058 210986 536294
rect 211222 536058 211306 536294
rect 211542 536058 211574 536294
rect 210954 509939 211574 536058
rect 217794 704838 218414 705830
rect 217794 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 218414 704838
rect 217794 704518 218414 704602
rect 217794 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 218414 704518
rect 217794 687454 218414 704282
rect 217794 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 218414 687454
rect 217794 687134 218414 687218
rect 217794 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 218414 687134
rect 217794 651454 218414 686898
rect 217794 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 218414 651454
rect 217794 651134 218414 651218
rect 217794 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 218414 651134
rect 217794 615454 218414 650898
rect 217794 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 218414 615454
rect 217794 615134 218414 615218
rect 217794 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 218414 615134
rect 217794 579454 218414 614898
rect 217794 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 218414 579454
rect 217794 579134 218414 579218
rect 217794 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 218414 579134
rect 217794 543454 218414 578898
rect 217794 543218 217826 543454
rect 218062 543218 218146 543454
rect 218382 543218 218414 543454
rect 217794 543134 218414 543218
rect 217794 542898 217826 543134
rect 218062 542898 218146 543134
rect 218382 542898 218414 543134
rect 217794 509939 218414 542898
rect 221514 691174 222134 706202
rect 221514 690938 221546 691174
rect 221782 690938 221866 691174
rect 222102 690938 222134 691174
rect 221514 690854 222134 690938
rect 221514 690618 221546 690854
rect 221782 690618 221866 690854
rect 222102 690618 222134 690854
rect 221514 655174 222134 690618
rect 221514 654938 221546 655174
rect 221782 654938 221866 655174
rect 222102 654938 222134 655174
rect 221514 654854 222134 654938
rect 221514 654618 221546 654854
rect 221782 654618 221866 654854
rect 222102 654618 222134 654854
rect 221514 619174 222134 654618
rect 221514 618938 221546 619174
rect 221782 618938 221866 619174
rect 222102 618938 222134 619174
rect 221514 618854 222134 618938
rect 221514 618618 221546 618854
rect 221782 618618 221866 618854
rect 222102 618618 222134 618854
rect 221514 583174 222134 618618
rect 221514 582938 221546 583174
rect 221782 582938 221866 583174
rect 222102 582938 222134 583174
rect 221514 582854 222134 582938
rect 221514 582618 221546 582854
rect 221782 582618 221866 582854
rect 222102 582618 222134 582854
rect 221514 547174 222134 582618
rect 221514 546938 221546 547174
rect 221782 546938 221866 547174
rect 222102 546938 222134 547174
rect 221514 546854 222134 546938
rect 221514 546618 221546 546854
rect 221782 546618 221866 546854
rect 222102 546618 222134 546854
rect 221514 511174 222134 546618
rect 221514 510938 221546 511174
rect 221782 510938 221866 511174
rect 222102 510938 222134 511174
rect 221514 510854 222134 510938
rect 221514 510618 221546 510854
rect 221782 510618 221866 510854
rect 222102 510618 222134 510854
rect 221514 509939 222134 510618
rect 225234 694894 225854 708122
rect 225234 694658 225266 694894
rect 225502 694658 225586 694894
rect 225822 694658 225854 694894
rect 225234 694574 225854 694658
rect 225234 694338 225266 694574
rect 225502 694338 225586 694574
rect 225822 694338 225854 694574
rect 225234 658894 225854 694338
rect 225234 658658 225266 658894
rect 225502 658658 225586 658894
rect 225822 658658 225854 658894
rect 225234 658574 225854 658658
rect 225234 658338 225266 658574
rect 225502 658338 225586 658574
rect 225822 658338 225854 658574
rect 225234 622894 225854 658338
rect 225234 622658 225266 622894
rect 225502 622658 225586 622894
rect 225822 622658 225854 622894
rect 225234 622574 225854 622658
rect 225234 622338 225266 622574
rect 225502 622338 225586 622574
rect 225822 622338 225854 622574
rect 225234 586894 225854 622338
rect 225234 586658 225266 586894
rect 225502 586658 225586 586894
rect 225822 586658 225854 586894
rect 225234 586574 225854 586658
rect 225234 586338 225266 586574
rect 225502 586338 225586 586574
rect 225822 586338 225854 586574
rect 225234 550894 225854 586338
rect 225234 550658 225266 550894
rect 225502 550658 225586 550894
rect 225822 550658 225854 550894
rect 225234 550574 225854 550658
rect 225234 550338 225266 550574
rect 225502 550338 225586 550574
rect 225822 550338 225854 550574
rect 225234 514894 225854 550338
rect 225234 514658 225266 514894
rect 225502 514658 225586 514894
rect 225822 514658 225854 514894
rect 225234 514574 225854 514658
rect 225234 514338 225266 514574
rect 225502 514338 225586 514574
rect 225822 514338 225854 514574
rect 225234 509939 225854 514338
rect 228954 698614 229574 710042
rect 246954 711558 247574 711590
rect 246954 711322 246986 711558
rect 247222 711322 247306 711558
rect 247542 711322 247574 711558
rect 246954 711238 247574 711322
rect 246954 711002 246986 711238
rect 247222 711002 247306 711238
rect 247542 711002 247574 711238
rect 243234 709638 243854 709670
rect 243234 709402 243266 709638
rect 243502 709402 243586 709638
rect 243822 709402 243854 709638
rect 243234 709318 243854 709402
rect 243234 709082 243266 709318
rect 243502 709082 243586 709318
rect 243822 709082 243854 709318
rect 239514 707718 240134 707750
rect 239514 707482 239546 707718
rect 239782 707482 239866 707718
rect 240102 707482 240134 707718
rect 239514 707398 240134 707482
rect 239514 707162 239546 707398
rect 239782 707162 239866 707398
rect 240102 707162 240134 707398
rect 228954 698378 228986 698614
rect 229222 698378 229306 698614
rect 229542 698378 229574 698614
rect 228954 698294 229574 698378
rect 228954 698058 228986 698294
rect 229222 698058 229306 698294
rect 229542 698058 229574 698294
rect 228954 662614 229574 698058
rect 228954 662378 228986 662614
rect 229222 662378 229306 662614
rect 229542 662378 229574 662614
rect 228954 662294 229574 662378
rect 228954 662058 228986 662294
rect 229222 662058 229306 662294
rect 229542 662058 229574 662294
rect 228954 626614 229574 662058
rect 228954 626378 228986 626614
rect 229222 626378 229306 626614
rect 229542 626378 229574 626614
rect 228954 626294 229574 626378
rect 228954 626058 228986 626294
rect 229222 626058 229306 626294
rect 229542 626058 229574 626294
rect 228954 590614 229574 626058
rect 228954 590378 228986 590614
rect 229222 590378 229306 590614
rect 229542 590378 229574 590614
rect 228954 590294 229574 590378
rect 228954 590058 228986 590294
rect 229222 590058 229306 590294
rect 229542 590058 229574 590294
rect 228954 554614 229574 590058
rect 228954 554378 228986 554614
rect 229222 554378 229306 554614
rect 229542 554378 229574 554614
rect 228954 554294 229574 554378
rect 228954 554058 228986 554294
rect 229222 554058 229306 554294
rect 229542 554058 229574 554294
rect 228954 518614 229574 554058
rect 228954 518378 228986 518614
rect 229222 518378 229306 518614
rect 229542 518378 229574 518614
rect 228954 518294 229574 518378
rect 228954 518058 228986 518294
rect 229222 518058 229306 518294
rect 229542 518058 229574 518294
rect 228954 509939 229574 518058
rect 235794 705798 236414 705830
rect 235794 705562 235826 705798
rect 236062 705562 236146 705798
rect 236382 705562 236414 705798
rect 235794 705478 236414 705562
rect 235794 705242 235826 705478
rect 236062 705242 236146 705478
rect 236382 705242 236414 705478
rect 235794 669454 236414 705242
rect 235794 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 236414 669454
rect 235794 669134 236414 669218
rect 235794 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 236414 669134
rect 235794 633454 236414 668898
rect 235794 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 236414 633454
rect 235794 633134 236414 633218
rect 235794 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 236414 633134
rect 235794 597454 236414 632898
rect 235794 597218 235826 597454
rect 236062 597218 236146 597454
rect 236382 597218 236414 597454
rect 235794 597134 236414 597218
rect 235794 596898 235826 597134
rect 236062 596898 236146 597134
rect 236382 596898 236414 597134
rect 235794 561454 236414 596898
rect 235794 561218 235826 561454
rect 236062 561218 236146 561454
rect 236382 561218 236414 561454
rect 235794 561134 236414 561218
rect 235794 560898 235826 561134
rect 236062 560898 236146 561134
rect 236382 560898 236414 561134
rect 235794 525454 236414 560898
rect 235794 525218 235826 525454
rect 236062 525218 236146 525454
rect 236382 525218 236414 525454
rect 235794 525134 236414 525218
rect 235794 524898 235826 525134
rect 236062 524898 236146 525134
rect 236382 524898 236414 525134
rect 235794 509939 236414 524898
rect 239514 673174 240134 707162
rect 239514 672938 239546 673174
rect 239782 672938 239866 673174
rect 240102 672938 240134 673174
rect 239514 672854 240134 672938
rect 239514 672618 239546 672854
rect 239782 672618 239866 672854
rect 240102 672618 240134 672854
rect 239514 637174 240134 672618
rect 239514 636938 239546 637174
rect 239782 636938 239866 637174
rect 240102 636938 240134 637174
rect 239514 636854 240134 636938
rect 239514 636618 239546 636854
rect 239782 636618 239866 636854
rect 240102 636618 240134 636854
rect 239514 601174 240134 636618
rect 239514 600938 239546 601174
rect 239782 600938 239866 601174
rect 240102 600938 240134 601174
rect 239514 600854 240134 600938
rect 239514 600618 239546 600854
rect 239782 600618 239866 600854
rect 240102 600618 240134 600854
rect 239514 565174 240134 600618
rect 239514 564938 239546 565174
rect 239782 564938 239866 565174
rect 240102 564938 240134 565174
rect 239514 564854 240134 564938
rect 239514 564618 239546 564854
rect 239782 564618 239866 564854
rect 240102 564618 240134 564854
rect 239514 529174 240134 564618
rect 239514 528938 239546 529174
rect 239782 528938 239866 529174
rect 240102 528938 240134 529174
rect 239514 528854 240134 528938
rect 239514 528618 239546 528854
rect 239782 528618 239866 528854
rect 240102 528618 240134 528854
rect 239514 509939 240134 528618
rect 243234 676894 243854 709082
rect 243234 676658 243266 676894
rect 243502 676658 243586 676894
rect 243822 676658 243854 676894
rect 243234 676574 243854 676658
rect 243234 676338 243266 676574
rect 243502 676338 243586 676574
rect 243822 676338 243854 676574
rect 243234 640894 243854 676338
rect 243234 640658 243266 640894
rect 243502 640658 243586 640894
rect 243822 640658 243854 640894
rect 243234 640574 243854 640658
rect 243234 640338 243266 640574
rect 243502 640338 243586 640574
rect 243822 640338 243854 640574
rect 243234 604894 243854 640338
rect 243234 604658 243266 604894
rect 243502 604658 243586 604894
rect 243822 604658 243854 604894
rect 243234 604574 243854 604658
rect 243234 604338 243266 604574
rect 243502 604338 243586 604574
rect 243822 604338 243854 604574
rect 243234 568894 243854 604338
rect 243234 568658 243266 568894
rect 243502 568658 243586 568894
rect 243822 568658 243854 568894
rect 243234 568574 243854 568658
rect 243234 568338 243266 568574
rect 243502 568338 243586 568574
rect 243822 568338 243854 568574
rect 243234 532894 243854 568338
rect 243234 532658 243266 532894
rect 243502 532658 243586 532894
rect 243822 532658 243854 532894
rect 243234 532574 243854 532658
rect 243234 532338 243266 532574
rect 243502 532338 243586 532574
rect 243822 532338 243854 532574
rect 243234 509939 243854 532338
rect 246954 680614 247574 711002
rect 264954 710598 265574 711590
rect 264954 710362 264986 710598
rect 265222 710362 265306 710598
rect 265542 710362 265574 710598
rect 264954 710278 265574 710362
rect 264954 710042 264986 710278
rect 265222 710042 265306 710278
rect 265542 710042 265574 710278
rect 261234 708678 261854 709670
rect 261234 708442 261266 708678
rect 261502 708442 261586 708678
rect 261822 708442 261854 708678
rect 261234 708358 261854 708442
rect 261234 708122 261266 708358
rect 261502 708122 261586 708358
rect 261822 708122 261854 708358
rect 257514 706758 258134 707750
rect 257514 706522 257546 706758
rect 257782 706522 257866 706758
rect 258102 706522 258134 706758
rect 257514 706438 258134 706522
rect 257514 706202 257546 706438
rect 257782 706202 257866 706438
rect 258102 706202 258134 706438
rect 246954 680378 246986 680614
rect 247222 680378 247306 680614
rect 247542 680378 247574 680614
rect 246954 680294 247574 680378
rect 246954 680058 246986 680294
rect 247222 680058 247306 680294
rect 247542 680058 247574 680294
rect 246954 644614 247574 680058
rect 246954 644378 246986 644614
rect 247222 644378 247306 644614
rect 247542 644378 247574 644614
rect 246954 644294 247574 644378
rect 246954 644058 246986 644294
rect 247222 644058 247306 644294
rect 247542 644058 247574 644294
rect 246954 608614 247574 644058
rect 246954 608378 246986 608614
rect 247222 608378 247306 608614
rect 247542 608378 247574 608614
rect 246954 608294 247574 608378
rect 246954 608058 246986 608294
rect 247222 608058 247306 608294
rect 247542 608058 247574 608294
rect 246954 572614 247574 608058
rect 246954 572378 246986 572614
rect 247222 572378 247306 572614
rect 247542 572378 247574 572614
rect 246954 572294 247574 572378
rect 246954 572058 246986 572294
rect 247222 572058 247306 572294
rect 247542 572058 247574 572294
rect 246954 536614 247574 572058
rect 246954 536378 246986 536614
rect 247222 536378 247306 536614
rect 247542 536378 247574 536614
rect 246954 536294 247574 536378
rect 246954 536058 246986 536294
rect 247222 536058 247306 536294
rect 247542 536058 247574 536294
rect 246954 509939 247574 536058
rect 253794 704838 254414 705830
rect 253794 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 254414 704838
rect 253794 704518 254414 704602
rect 253794 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 254414 704518
rect 253794 687454 254414 704282
rect 253794 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 254414 687454
rect 253794 687134 254414 687218
rect 253794 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 254414 687134
rect 253794 651454 254414 686898
rect 253794 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 254414 651454
rect 253794 651134 254414 651218
rect 253794 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 254414 651134
rect 253794 615454 254414 650898
rect 253794 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 254414 615454
rect 253794 615134 254414 615218
rect 253794 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 254414 615134
rect 253794 579454 254414 614898
rect 253794 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 254414 579454
rect 253794 579134 254414 579218
rect 253794 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 254414 579134
rect 253794 543454 254414 578898
rect 253794 543218 253826 543454
rect 254062 543218 254146 543454
rect 254382 543218 254414 543454
rect 253794 543134 254414 543218
rect 253794 542898 253826 543134
rect 254062 542898 254146 543134
rect 254382 542898 254414 543134
rect 253794 509939 254414 542898
rect 257514 691174 258134 706202
rect 257514 690938 257546 691174
rect 257782 690938 257866 691174
rect 258102 690938 258134 691174
rect 257514 690854 258134 690938
rect 257514 690618 257546 690854
rect 257782 690618 257866 690854
rect 258102 690618 258134 690854
rect 257514 655174 258134 690618
rect 257514 654938 257546 655174
rect 257782 654938 257866 655174
rect 258102 654938 258134 655174
rect 257514 654854 258134 654938
rect 257514 654618 257546 654854
rect 257782 654618 257866 654854
rect 258102 654618 258134 654854
rect 257514 619174 258134 654618
rect 257514 618938 257546 619174
rect 257782 618938 257866 619174
rect 258102 618938 258134 619174
rect 257514 618854 258134 618938
rect 257514 618618 257546 618854
rect 257782 618618 257866 618854
rect 258102 618618 258134 618854
rect 257514 583174 258134 618618
rect 257514 582938 257546 583174
rect 257782 582938 257866 583174
rect 258102 582938 258134 583174
rect 257514 582854 258134 582938
rect 257514 582618 257546 582854
rect 257782 582618 257866 582854
rect 258102 582618 258134 582854
rect 257514 547174 258134 582618
rect 257514 546938 257546 547174
rect 257782 546938 257866 547174
rect 258102 546938 258134 547174
rect 257514 546854 258134 546938
rect 257514 546618 257546 546854
rect 257782 546618 257866 546854
rect 258102 546618 258134 546854
rect 257514 511174 258134 546618
rect 257514 510938 257546 511174
rect 257782 510938 257866 511174
rect 258102 510938 258134 511174
rect 257514 510854 258134 510938
rect 257514 510618 257546 510854
rect 257782 510618 257866 510854
rect 258102 510618 258134 510854
rect 257514 509939 258134 510618
rect 261234 694894 261854 708122
rect 261234 694658 261266 694894
rect 261502 694658 261586 694894
rect 261822 694658 261854 694894
rect 261234 694574 261854 694658
rect 261234 694338 261266 694574
rect 261502 694338 261586 694574
rect 261822 694338 261854 694574
rect 261234 658894 261854 694338
rect 261234 658658 261266 658894
rect 261502 658658 261586 658894
rect 261822 658658 261854 658894
rect 261234 658574 261854 658658
rect 261234 658338 261266 658574
rect 261502 658338 261586 658574
rect 261822 658338 261854 658574
rect 261234 622894 261854 658338
rect 261234 622658 261266 622894
rect 261502 622658 261586 622894
rect 261822 622658 261854 622894
rect 261234 622574 261854 622658
rect 261234 622338 261266 622574
rect 261502 622338 261586 622574
rect 261822 622338 261854 622574
rect 261234 586894 261854 622338
rect 261234 586658 261266 586894
rect 261502 586658 261586 586894
rect 261822 586658 261854 586894
rect 261234 586574 261854 586658
rect 261234 586338 261266 586574
rect 261502 586338 261586 586574
rect 261822 586338 261854 586574
rect 261234 550894 261854 586338
rect 261234 550658 261266 550894
rect 261502 550658 261586 550894
rect 261822 550658 261854 550894
rect 261234 550574 261854 550658
rect 261234 550338 261266 550574
rect 261502 550338 261586 550574
rect 261822 550338 261854 550574
rect 261234 514894 261854 550338
rect 261234 514658 261266 514894
rect 261502 514658 261586 514894
rect 261822 514658 261854 514894
rect 261234 514574 261854 514658
rect 261234 514338 261266 514574
rect 261502 514338 261586 514574
rect 261822 514338 261854 514574
rect 261234 509939 261854 514338
rect 264954 698614 265574 710042
rect 282954 711558 283574 711590
rect 282954 711322 282986 711558
rect 283222 711322 283306 711558
rect 283542 711322 283574 711558
rect 282954 711238 283574 711322
rect 282954 711002 282986 711238
rect 283222 711002 283306 711238
rect 283542 711002 283574 711238
rect 279234 709638 279854 709670
rect 279234 709402 279266 709638
rect 279502 709402 279586 709638
rect 279822 709402 279854 709638
rect 279234 709318 279854 709402
rect 279234 709082 279266 709318
rect 279502 709082 279586 709318
rect 279822 709082 279854 709318
rect 275514 707718 276134 707750
rect 275514 707482 275546 707718
rect 275782 707482 275866 707718
rect 276102 707482 276134 707718
rect 275514 707398 276134 707482
rect 275514 707162 275546 707398
rect 275782 707162 275866 707398
rect 276102 707162 276134 707398
rect 264954 698378 264986 698614
rect 265222 698378 265306 698614
rect 265542 698378 265574 698614
rect 264954 698294 265574 698378
rect 264954 698058 264986 698294
rect 265222 698058 265306 698294
rect 265542 698058 265574 698294
rect 264954 662614 265574 698058
rect 264954 662378 264986 662614
rect 265222 662378 265306 662614
rect 265542 662378 265574 662614
rect 264954 662294 265574 662378
rect 264954 662058 264986 662294
rect 265222 662058 265306 662294
rect 265542 662058 265574 662294
rect 264954 626614 265574 662058
rect 264954 626378 264986 626614
rect 265222 626378 265306 626614
rect 265542 626378 265574 626614
rect 264954 626294 265574 626378
rect 264954 626058 264986 626294
rect 265222 626058 265306 626294
rect 265542 626058 265574 626294
rect 264954 590614 265574 626058
rect 264954 590378 264986 590614
rect 265222 590378 265306 590614
rect 265542 590378 265574 590614
rect 264954 590294 265574 590378
rect 264954 590058 264986 590294
rect 265222 590058 265306 590294
rect 265542 590058 265574 590294
rect 264954 554614 265574 590058
rect 264954 554378 264986 554614
rect 265222 554378 265306 554614
rect 265542 554378 265574 554614
rect 264954 554294 265574 554378
rect 264954 554058 264986 554294
rect 265222 554058 265306 554294
rect 265542 554058 265574 554294
rect 264954 518614 265574 554058
rect 264954 518378 264986 518614
rect 265222 518378 265306 518614
rect 265542 518378 265574 518614
rect 264954 518294 265574 518378
rect 264954 518058 264986 518294
rect 265222 518058 265306 518294
rect 265542 518058 265574 518294
rect 264954 509939 265574 518058
rect 271794 705798 272414 705830
rect 271794 705562 271826 705798
rect 272062 705562 272146 705798
rect 272382 705562 272414 705798
rect 271794 705478 272414 705562
rect 271794 705242 271826 705478
rect 272062 705242 272146 705478
rect 272382 705242 272414 705478
rect 271794 669454 272414 705242
rect 271794 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 272414 669454
rect 271794 669134 272414 669218
rect 271794 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 272414 669134
rect 271794 633454 272414 668898
rect 271794 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 272414 633454
rect 271794 633134 272414 633218
rect 271794 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 272414 633134
rect 271794 597454 272414 632898
rect 271794 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 272414 597454
rect 271794 597134 272414 597218
rect 271794 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 272414 597134
rect 271794 561454 272414 596898
rect 271794 561218 271826 561454
rect 272062 561218 272146 561454
rect 272382 561218 272414 561454
rect 271794 561134 272414 561218
rect 271794 560898 271826 561134
rect 272062 560898 272146 561134
rect 272382 560898 272414 561134
rect 271794 525454 272414 560898
rect 271794 525218 271826 525454
rect 272062 525218 272146 525454
rect 272382 525218 272414 525454
rect 271794 525134 272414 525218
rect 271794 524898 271826 525134
rect 272062 524898 272146 525134
rect 272382 524898 272414 525134
rect 271794 509939 272414 524898
rect 275514 673174 276134 707162
rect 275514 672938 275546 673174
rect 275782 672938 275866 673174
rect 276102 672938 276134 673174
rect 275514 672854 276134 672938
rect 275514 672618 275546 672854
rect 275782 672618 275866 672854
rect 276102 672618 276134 672854
rect 275514 637174 276134 672618
rect 275514 636938 275546 637174
rect 275782 636938 275866 637174
rect 276102 636938 276134 637174
rect 275514 636854 276134 636938
rect 275514 636618 275546 636854
rect 275782 636618 275866 636854
rect 276102 636618 276134 636854
rect 275514 601174 276134 636618
rect 275514 600938 275546 601174
rect 275782 600938 275866 601174
rect 276102 600938 276134 601174
rect 275514 600854 276134 600938
rect 275514 600618 275546 600854
rect 275782 600618 275866 600854
rect 276102 600618 276134 600854
rect 275514 565174 276134 600618
rect 275514 564938 275546 565174
rect 275782 564938 275866 565174
rect 276102 564938 276134 565174
rect 275514 564854 276134 564938
rect 275514 564618 275546 564854
rect 275782 564618 275866 564854
rect 276102 564618 276134 564854
rect 275514 529174 276134 564618
rect 275514 528938 275546 529174
rect 275782 528938 275866 529174
rect 276102 528938 276134 529174
rect 275514 528854 276134 528938
rect 275514 528618 275546 528854
rect 275782 528618 275866 528854
rect 276102 528618 276134 528854
rect 275514 509939 276134 528618
rect 279234 676894 279854 709082
rect 279234 676658 279266 676894
rect 279502 676658 279586 676894
rect 279822 676658 279854 676894
rect 279234 676574 279854 676658
rect 279234 676338 279266 676574
rect 279502 676338 279586 676574
rect 279822 676338 279854 676574
rect 279234 640894 279854 676338
rect 279234 640658 279266 640894
rect 279502 640658 279586 640894
rect 279822 640658 279854 640894
rect 279234 640574 279854 640658
rect 279234 640338 279266 640574
rect 279502 640338 279586 640574
rect 279822 640338 279854 640574
rect 279234 604894 279854 640338
rect 279234 604658 279266 604894
rect 279502 604658 279586 604894
rect 279822 604658 279854 604894
rect 279234 604574 279854 604658
rect 279234 604338 279266 604574
rect 279502 604338 279586 604574
rect 279822 604338 279854 604574
rect 279234 568894 279854 604338
rect 279234 568658 279266 568894
rect 279502 568658 279586 568894
rect 279822 568658 279854 568894
rect 279234 568574 279854 568658
rect 279234 568338 279266 568574
rect 279502 568338 279586 568574
rect 279822 568338 279854 568574
rect 279234 532894 279854 568338
rect 279234 532658 279266 532894
rect 279502 532658 279586 532894
rect 279822 532658 279854 532894
rect 279234 532574 279854 532658
rect 279234 532338 279266 532574
rect 279502 532338 279586 532574
rect 279822 532338 279854 532574
rect 279234 509939 279854 532338
rect 282954 680614 283574 711002
rect 300954 710598 301574 711590
rect 300954 710362 300986 710598
rect 301222 710362 301306 710598
rect 301542 710362 301574 710598
rect 300954 710278 301574 710362
rect 300954 710042 300986 710278
rect 301222 710042 301306 710278
rect 301542 710042 301574 710278
rect 297234 708678 297854 709670
rect 297234 708442 297266 708678
rect 297502 708442 297586 708678
rect 297822 708442 297854 708678
rect 297234 708358 297854 708442
rect 297234 708122 297266 708358
rect 297502 708122 297586 708358
rect 297822 708122 297854 708358
rect 293514 706758 294134 707750
rect 293514 706522 293546 706758
rect 293782 706522 293866 706758
rect 294102 706522 294134 706758
rect 293514 706438 294134 706522
rect 293514 706202 293546 706438
rect 293782 706202 293866 706438
rect 294102 706202 294134 706438
rect 282954 680378 282986 680614
rect 283222 680378 283306 680614
rect 283542 680378 283574 680614
rect 282954 680294 283574 680378
rect 282954 680058 282986 680294
rect 283222 680058 283306 680294
rect 283542 680058 283574 680294
rect 282954 644614 283574 680058
rect 282954 644378 282986 644614
rect 283222 644378 283306 644614
rect 283542 644378 283574 644614
rect 282954 644294 283574 644378
rect 282954 644058 282986 644294
rect 283222 644058 283306 644294
rect 283542 644058 283574 644294
rect 282954 608614 283574 644058
rect 282954 608378 282986 608614
rect 283222 608378 283306 608614
rect 283542 608378 283574 608614
rect 282954 608294 283574 608378
rect 282954 608058 282986 608294
rect 283222 608058 283306 608294
rect 283542 608058 283574 608294
rect 282954 572614 283574 608058
rect 282954 572378 282986 572614
rect 283222 572378 283306 572614
rect 283542 572378 283574 572614
rect 282954 572294 283574 572378
rect 282954 572058 282986 572294
rect 283222 572058 283306 572294
rect 283542 572058 283574 572294
rect 282954 536614 283574 572058
rect 282954 536378 282986 536614
rect 283222 536378 283306 536614
rect 283542 536378 283574 536614
rect 282954 536294 283574 536378
rect 282954 536058 282986 536294
rect 283222 536058 283306 536294
rect 283542 536058 283574 536294
rect 282954 509939 283574 536058
rect 289794 704838 290414 705830
rect 289794 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 290414 704838
rect 289794 704518 290414 704602
rect 289794 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 290414 704518
rect 289794 687454 290414 704282
rect 289794 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 290414 687454
rect 289794 687134 290414 687218
rect 289794 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 290414 687134
rect 289794 651454 290414 686898
rect 289794 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 290414 651454
rect 289794 651134 290414 651218
rect 289794 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 290414 651134
rect 289794 615454 290414 650898
rect 289794 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 290414 615454
rect 289794 615134 290414 615218
rect 289794 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 290414 615134
rect 289794 579454 290414 614898
rect 289794 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 290414 579454
rect 289794 579134 290414 579218
rect 289794 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 290414 579134
rect 289794 543454 290414 578898
rect 289794 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 290414 543454
rect 289794 543134 290414 543218
rect 289794 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 290414 543134
rect 289794 509939 290414 542898
rect 293514 691174 294134 706202
rect 293514 690938 293546 691174
rect 293782 690938 293866 691174
rect 294102 690938 294134 691174
rect 293514 690854 294134 690938
rect 293514 690618 293546 690854
rect 293782 690618 293866 690854
rect 294102 690618 294134 690854
rect 293514 655174 294134 690618
rect 293514 654938 293546 655174
rect 293782 654938 293866 655174
rect 294102 654938 294134 655174
rect 293514 654854 294134 654938
rect 293514 654618 293546 654854
rect 293782 654618 293866 654854
rect 294102 654618 294134 654854
rect 293514 619174 294134 654618
rect 293514 618938 293546 619174
rect 293782 618938 293866 619174
rect 294102 618938 294134 619174
rect 293514 618854 294134 618938
rect 293514 618618 293546 618854
rect 293782 618618 293866 618854
rect 294102 618618 294134 618854
rect 293514 583174 294134 618618
rect 293514 582938 293546 583174
rect 293782 582938 293866 583174
rect 294102 582938 294134 583174
rect 293514 582854 294134 582938
rect 293514 582618 293546 582854
rect 293782 582618 293866 582854
rect 294102 582618 294134 582854
rect 293514 547174 294134 582618
rect 293514 546938 293546 547174
rect 293782 546938 293866 547174
rect 294102 546938 294134 547174
rect 293514 546854 294134 546938
rect 293514 546618 293546 546854
rect 293782 546618 293866 546854
rect 294102 546618 294134 546854
rect 293514 511174 294134 546618
rect 293514 510938 293546 511174
rect 293782 510938 293866 511174
rect 294102 510938 294134 511174
rect 293514 510854 294134 510938
rect 293514 510618 293546 510854
rect 293782 510618 293866 510854
rect 294102 510618 294134 510854
rect 293514 509939 294134 510618
rect 297234 694894 297854 708122
rect 297234 694658 297266 694894
rect 297502 694658 297586 694894
rect 297822 694658 297854 694894
rect 297234 694574 297854 694658
rect 297234 694338 297266 694574
rect 297502 694338 297586 694574
rect 297822 694338 297854 694574
rect 297234 658894 297854 694338
rect 297234 658658 297266 658894
rect 297502 658658 297586 658894
rect 297822 658658 297854 658894
rect 297234 658574 297854 658658
rect 297234 658338 297266 658574
rect 297502 658338 297586 658574
rect 297822 658338 297854 658574
rect 297234 622894 297854 658338
rect 297234 622658 297266 622894
rect 297502 622658 297586 622894
rect 297822 622658 297854 622894
rect 297234 622574 297854 622658
rect 297234 622338 297266 622574
rect 297502 622338 297586 622574
rect 297822 622338 297854 622574
rect 297234 586894 297854 622338
rect 297234 586658 297266 586894
rect 297502 586658 297586 586894
rect 297822 586658 297854 586894
rect 297234 586574 297854 586658
rect 297234 586338 297266 586574
rect 297502 586338 297586 586574
rect 297822 586338 297854 586574
rect 297234 550894 297854 586338
rect 297234 550658 297266 550894
rect 297502 550658 297586 550894
rect 297822 550658 297854 550894
rect 297234 550574 297854 550658
rect 297234 550338 297266 550574
rect 297502 550338 297586 550574
rect 297822 550338 297854 550574
rect 297234 514894 297854 550338
rect 297234 514658 297266 514894
rect 297502 514658 297586 514894
rect 297822 514658 297854 514894
rect 297234 514574 297854 514658
rect 297234 514338 297266 514574
rect 297502 514338 297586 514574
rect 297822 514338 297854 514574
rect 297234 509939 297854 514338
rect 300954 698614 301574 710042
rect 318954 711558 319574 711590
rect 318954 711322 318986 711558
rect 319222 711322 319306 711558
rect 319542 711322 319574 711558
rect 318954 711238 319574 711322
rect 318954 711002 318986 711238
rect 319222 711002 319306 711238
rect 319542 711002 319574 711238
rect 315234 709638 315854 709670
rect 315234 709402 315266 709638
rect 315502 709402 315586 709638
rect 315822 709402 315854 709638
rect 315234 709318 315854 709402
rect 315234 709082 315266 709318
rect 315502 709082 315586 709318
rect 315822 709082 315854 709318
rect 311514 707718 312134 707750
rect 311514 707482 311546 707718
rect 311782 707482 311866 707718
rect 312102 707482 312134 707718
rect 311514 707398 312134 707482
rect 311514 707162 311546 707398
rect 311782 707162 311866 707398
rect 312102 707162 312134 707398
rect 300954 698378 300986 698614
rect 301222 698378 301306 698614
rect 301542 698378 301574 698614
rect 300954 698294 301574 698378
rect 300954 698058 300986 698294
rect 301222 698058 301306 698294
rect 301542 698058 301574 698294
rect 300954 662614 301574 698058
rect 300954 662378 300986 662614
rect 301222 662378 301306 662614
rect 301542 662378 301574 662614
rect 300954 662294 301574 662378
rect 300954 662058 300986 662294
rect 301222 662058 301306 662294
rect 301542 662058 301574 662294
rect 300954 626614 301574 662058
rect 300954 626378 300986 626614
rect 301222 626378 301306 626614
rect 301542 626378 301574 626614
rect 300954 626294 301574 626378
rect 300954 626058 300986 626294
rect 301222 626058 301306 626294
rect 301542 626058 301574 626294
rect 300954 590614 301574 626058
rect 300954 590378 300986 590614
rect 301222 590378 301306 590614
rect 301542 590378 301574 590614
rect 300954 590294 301574 590378
rect 300954 590058 300986 590294
rect 301222 590058 301306 590294
rect 301542 590058 301574 590294
rect 300954 554614 301574 590058
rect 300954 554378 300986 554614
rect 301222 554378 301306 554614
rect 301542 554378 301574 554614
rect 300954 554294 301574 554378
rect 300954 554058 300986 554294
rect 301222 554058 301306 554294
rect 301542 554058 301574 554294
rect 300954 518614 301574 554058
rect 300954 518378 300986 518614
rect 301222 518378 301306 518614
rect 301542 518378 301574 518614
rect 300954 518294 301574 518378
rect 300954 518058 300986 518294
rect 301222 518058 301306 518294
rect 301542 518058 301574 518294
rect 300954 509939 301574 518058
rect 307794 705798 308414 705830
rect 307794 705562 307826 705798
rect 308062 705562 308146 705798
rect 308382 705562 308414 705798
rect 307794 705478 308414 705562
rect 307794 705242 307826 705478
rect 308062 705242 308146 705478
rect 308382 705242 308414 705478
rect 307794 669454 308414 705242
rect 307794 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 308414 669454
rect 307794 669134 308414 669218
rect 307794 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 308414 669134
rect 307794 633454 308414 668898
rect 307794 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 308414 633454
rect 307794 633134 308414 633218
rect 307794 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 308414 633134
rect 307794 597454 308414 632898
rect 307794 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 308414 597454
rect 307794 597134 308414 597218
rect 307794 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 308414 597134
rect 307794 561454 308414 596898
rect 307794 561218 307826 561454
rect 308062 561218 308146 561454
rect 308382 561218 308414 561454
rect 307794 561134 308414 561218
rect 307794 560898 307826 561134
rect 308062 560898 308146 561134
rect 308382 560898 308414 561134
rect 307794 525454 308414 560898
rect 307794 525218 307826 525454
rect 308062 525218 308146 525454
rect 308382 525218 308414 525454
rect 307794 525134 308414 525218
rect 307794 524898 307826 525134
rect 308062 524898 308146 525134
rect 308382 524898 308414 525134
rect 307794 509939 308414 524898
rect 311514 673174 312134 707162
rect 311514 672938 311546 673174
rect 311782 672938 311866 673174
rect 312102 672938 312134 673174
rect 311514 672854 312134 672938
rect 311514 672618 311546 672854
rect 311782 672618 311866 672854
rect 312102 672618 312134 672854
rect 311514 637174 312134 672618
rect 311514 636938 311546 637174
rect 311782 636938 311866 637174
rect 312102 636938 312134 637174
rect 311514 636854 312134 636938
rect 311514 636618 311546 636854
rect 311782 636618 311866 636854
rect 312102 636618 312134 636854
rect 311514 601174 312134 636618
rect 311514 600938 311546 601174
rect 311782 600938 311866 601174
rect 312102 600938 312134 601174
rect 311514 600854 312134 600938
rect 311514 600618 311546 600854
rect 311782 600618 311866 600854
rect 312102 600618 312134 600854
rect 311514 565174 312134 600618
rect 311514 564938 311546 565174
rect 311782 564938 311866 565174
rect 312102 564938 312134 565174
rect 311514 564854 312134 564938
rect 311514 564618 311546 564854
rect 311782 564618 311866 564854
rect 312102 564618 312134 564854
rect 311514 529174 312134 564618
rect 311514 528938 311546 529174
rect 311782 528938 311866 529174
rect 312102 528938 312134 529174
rect 311514 528854 312134 528938
rect 311514 528618 311546 528854
rect 311782 528618 311866 528854
rect 312102 528618 312134 528854
rect 311514 509939 312134 528618
rect 315234 676894 315854 709082
rect 315234 676658 315266 676894
rect 315502 676658 315586 676894
rect 315822 676658 315854 676894
rect 315234 676574 315854 676658
rect 315234 676338 315266 676574
rect 315502 676338 315586 676574
rect 315822 676338 315854 676574
rect 315234 640894 315854 676338
rect 315234 640658 315266 640894
rect 315502 640658 315586 640894
rect 315822 640658 315854 640894
rect 315234 640574 315854 640658
rect 315234 640338 315266 640574
rect 315502 640338 315586 640574
rect 315822 640338 315854 640574
rect 315234 604894 315854 640338
rect 315234 604658 315266 604894
rect 315502 604658 315586 604894
rect 315822 604658 315854 604894
rect 315234 604574 315854 604658
rect 315234 604338 315266 604574
rect 315502 604338 315586 604574
rect 315822 604338 315854 604574
rect 315234 568894 315854 604338
rect 315234 568658 315266 568894
rect 315502 568658 315586 568894
rect 315822 568658 315854 568894
rect 315234 568574 315854 568658
rect 315234 568338 315266 568574
rect 315502 568338 315586 568574
rect 315822 568338 315854 568574
rect 315234 532894 315854 568338
rect 315234 532658 315266 532894
rect 315502 532658 315586 532894
rect 315822 532658 315854 532894
rect 315234 532574 315854 532658
rect 315234 532338 315266 532574
rect 315502 532338 315586 532574
rect 315822 532338 315854 532574
rect 315234 509939 315854 532338
rect 318954 680614 319574 711002
rect 336954 710598 337574 711590
rect 336954 710362 336986 710598
rect 337222 710362 337306 710598
rect 337542 710362 337574 710598
rect 336954 710278 337574 710362
rect 336954 710042 336986 710278
rect 337222 710042 337306 710278
rect 337542 710042 337574 710278
rect 333234 708678 333854 709670
rect 333234 708442 333266 708678
rect 333502 708442 333586 708678
rect 333822 708442 333854 708678
rect 333234 708358 333854 708442
rect 333234 708122 333266 708358
rect 333502 708122 333586 708358
rect 333822 708122 333854 708358
rect 329514 706758 330134 707750
rect 329514 706522 329546 706758
rect 329782 706522 329866 706758
rect 330102 706522 330134 706758
rect 329514 706438 330134 706522
rect 329514 706202 329546 706438
rect 329782 706202 329866 706438
rect 330102 706202 330134 706438
rect 318954 680378 318986 680614
rect 319222 680378 319306 680614
rect 319542 680378 319574 680614
rect 318954 680294 319574 680378
rect 318954 680058 318986 680294
rect 319222 680058 319306 680294
rect 319542 680058 319574 680294
rect 318954 644614 319574 680058
rect 318954 644378 318986 644614
rect 319222 644378 319306 644614
rect 319542 644378 319574 644614
rect 318954 644294 319574 644378
rect 318954 644058 318986 644294
rect 319222 644058 319306 644294
rect 319542 644058 319574 644294
rect 318954 608614 319574 644058
rect 318954 608378 318986 608614
rect 319222 608378 319306 608614
rect 319542 608378 319574 608614
rect 318954 608294 319574 608378
rect 318954 608058 318986 608294
rect 319222 608058 319306 608294
rect 319542 608058 319574 608294
rect 318954 572614 319574 608058
rect 318954 572378 318986 572614
rect 319222 572378 319306 572614
rect 319542 572378 319574 572614
rect 318954 572294 319574 572378
rect 318954 572058 318986 572294
rect 319222 572058 319306 572294
rect 319542 572058 319574 572294
rect 318954 536614 319574 572058
rect 318954 536378 318986 536614
rect 319222 536378 319306 536614
rect 319542 536378 319574 536614
rect 318954 536294 319574 536378
rect 318954 536058 318986 536294
rect 319222 536058 319306 536294
rect 319542 536058 319574 536294
rect 318954 509939 319574 536058
rect 325794 704838 326414 705830
rect 325794 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 326414 704838
rect 325794 704518 326414 704602
rect 325794 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 326414 704518
rect 325794 687454 326414 704282
rect 325794 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 326414 687454
rect 325794 687134 326414 687218
rect 325794 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 326414 687134
rect 325794 651454 326414 686898
rect 325794 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 326414 651454
rect 325794 651134 326414 651218
rect 325794 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 326414 651134
rect 325794 615454 326414 650898
rect 325794 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 326414 615454
rect 325794 615134 326414 615218
rect 325794 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 326414 615134
rect 325794 579454 326414 614898
rect 325794 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 326414 579454
rect 325794 579134 326414 579218
rect 325794 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 326414 579134
rect 325794 543454 326414 578898
rect 325794 543218 325826 543454
rect 326062 543218 326146 543454
rect 326382 543218 326414 543454
rect 325794 543134 326414 543218
rect 325794 542898 325826 543134
rect 326062 542898 326146 543134
rect 326382 542898 326414 543134
rect 325794 509939 326414 542898
rect 329514 691174 330134 706202
rect 329514 690938 329546 691174
rect 329782 690938 329866 691174
rect 330102 690938 330134 691174
rect 329514 690854 330134 690938
rect 329514 690618 329546 690854
rect 329782 690618 329866 690854
rect 330102 690618 330134 690854
rect 329514 655174 330134 690618
rect 329514 654938 329546 655174
rect 329782 654938 329866 655174
rect 330102 654938 330134 655174
rect 329514 654854 330134 654938
rect 329514 654618 329546 654854
rect 329782 654618 329866 654854
rect 330102 654618 330134 654854
rect 329514 619174 330134 654618
rect 329514 618938 329546 619174
rect 329782 618938 329866 619174
rect 330102 618938 330134 619174
rect 329514 618854 330134 618938
rect 329514 618618 329546 618854
rect 329782 618618 329866 618854
rect 330102 618618 330134 618854
rect 329514 583174 330134 618618
rect 329514 582938 329546 583174
rect 329782 582938 329866 583174
rect 330102 582938 330134 583174
rect 329514 582854 330134 582938
rect 329514 582618 329546 582854
rect 329782 582618 329866 582854
rect 330102 582618 330134 582854
rect 329514 547174 330134 582618
rect 329514 546938 329546 547174
rect 329782 546938 329866 547174
rect 330102 546938 330134 547174
rect 329514 546854 330134 546938
rect 329514 546618 329546 546854
rect 329782 546618 329866 546854
rect 330102 546618 330134 546854
rect 329514 511174 330134 546618
rect 329514 510938 329546 511174
rect 329782 510938 329866 511174
rect 330102 510938 330134 511174
rect 329514 510854 330134 510938
rect 329514 510618 329546 510854
rect 329782 510618 329866 510854
rect 330102 510618 330134 510854
rect 329514 509939 330134 510618
rect 333234 694894 333854 708122
rect 333234 694658 333266 694894
rect 333502 694658 333586 694894
rect 333822 694658 333854 694894
rect 333234 694574 333854 694658
rect 333234 694338 333266 694574
rect 333502 694338 333586 694574
rect 333822 694338 333854 694574
rect 333234 658894 333854 694338
rect 333234 658658 333266 658894
rect 333502 658658 333586 658894
rect 333822 658658 333854 658894
rect 333234 658574 333854 658658
rect 333234 658338 333266 658574
rect 333502 658338 333586 658574
rect 333822 658338 333854 658574
rect 333234 622894 333854 658338
rect 333234 622658 333266 622894
rect 333502 622658 333586 622894
rect 333822 622658 333854 622894
rect 333234 622574 333854 622658
rect 333234 622338 333266 622574
rect 333502 622338 333586 622574
rect 333822 622338 333854 622574
rect 333234 586894 333854 622338
rect 333234 586658 333266 586894
rect 333502 586658 333586 586894
rect 333822 586658 333854 586894
rect 333234 586574 333854 586658
rect 333234 586338 333266 586574
rect 333502 586338 333586 586574
rect 333822 586338 333854 586574
rect 333234 550894 333854 586338
rect 333234 550658 333266 550894
rect 333502 550658 333586 550894
rect 333822 550658 333854 550894
rect 333234 550574 333854 550658
rect 333234 550338 333266 550574
rect 333502 550338 333586 550574
rect 333822 550338 333854 550574
rect 333234 514894 333854 550338
rect 333234 514658 333266 514894
rect 333502 514658 333586 514894
rect 333822 514658 333854 514894
rect 333234 514574 333854 514658
rect 333234 514338 333266 514574
rect 333502 514338 333586 514574
rect 333822 514338 333854 514574
rect 333234 509939 333854 514338
rect 336954 698614 337574 710042
rect 354954 711558 355574 711590
rect 354954 711322 354986 711558
rect 355222 711322 355306 711558
rect 355542 711322 355574 711558
rect 354954 711238 355574 711322
rect 354954 711002 354986 711238
rect 355222 711002 355306 711238
rect 355542 711002 355574 711238
rect 351234 709638 351854 709670
rect 351234 709402 351266 709638
rect 351502 709402 351586 709638
rect 351822 709402 351854 709638
rect 351234 709318 351854 709402
rect 351234 709082 351266 709318
rect 351502 709082 351586 709318
rect 351822 709082 351854 709318
rect 347514 707718 348134 707750
rect 347514 707482 347546 707718
rect 347782 707482 347866 707718
rect 348102 707482 348134 707718
rect 347514 707398 348134 707482
rect 347514 707162 347546 707398
rect 347782 707162 347866 707398
rect 348102 707162 348134 707398
rect 336954 698378 336986 698614
rect 337222 698378 337306 698614
rect 337542 698378 337574 698614
rect 336954 698294 337574 698378
rect 336954 698058 336986 698294
rect 337222 698058 337306 698294
rect 337542 698058 337574 698294
rect 336954 662614 337574 698058
rect 336954 662378 336986 662614
rect 337222 662378 337306 662614
rect 337542 662378 337574 662614
rect 336954 662294 337574 662378
rect 336954 662058 336986 662294
rect 337222 662058 337306 662294
rect 337542 662058 337574 662294
rect 336954 626614 337574 662058
rect 336954 626378 336986 626614
rect 337222 626378 337306 626614
rect 337542 626378 337574 626614
rect 336954 626294 337574 626378
rect 336954 626058 336986 626294
rect 337222 626058 337306 626294
rect 337542 626058 337574 626294
rect 336954 590614 337574 626058
rect 336954 590378 336986 590614
rect 337222 590378 337306 590614
rect 337542 590378 337574 590614
rect 336954 590294 337574 590378
rect 336954 590058 336986 590294
rect 337222 590058 337306 590294
rect 337542 590058 337574 590294
rect 336954 554614 337574 590058
rect 336954 554378 336986 554614
rect 337222 554378 337306 554614
rect 337542 554378 337574 554614
rect 336954 554294 337574 554378
rect 336954 554058 336986 554294
rect 337222 554058 337306 554294
rect 337542 554058 337574 554294
rect 336954 518614 337574 554058
rect 336954 518378 336986 518614
rect 337222 518378 337306 518614
rect 337542 518378 337574 518614
rect 336954 518294 337574 518378
rect 336954 518058 336986 518294
rect 337222 518058 337306 518294
rect 337542 518058 337574 518294
rect 336954 509939 337574 518058
rect 343794 705798 344414 705830
rect 343794 705562 343826 705798
rect 344062 705562 344146 705798
rect 344382 705562 344414 705798
rect 343794 705478 344414 705562
rect 343794 705242 343826 705478
rect 344062 705242 344146 705478
rect 344382 705242 344414 705478
rect 343794 669454 344414 705242
rect 343794 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 344414 669454
rect 343794 669134 344414 669218
rect 343794 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 344414 669134
rect 343794 633454 344414 668898
rect 343794 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 344414 633454
rect 343794 633134 344414 633218
rect 343794 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 344414 633134
rect 343794 597454 344414 632898
rect 343794 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 344414 597454
rect 343794 597134 344414 597218
rect 343794 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 344414 597134
rect 343794 561454 344414 596898
rect 343794 561218 343826 561454
rect 344062 561218 344146 561454
rect 344382 561218 344414 561454
rect 343794 561134 344414 561218
rect 343794 560898 343826 561134
rect 344062 560898 344146 561134
rect 344382 560898 344414 561134
rect 343794 525454 344414 560898
rect 343794 525218 343826 525454
rect 344062 525218 344146 525454
rect 344382 525218 344414 525454
rect 343794 525134 344414 525218
rect 343794 524898 343826 525134
rect 344062 524898 344146 525134
rect 344382 524898 344414 525134
rect 343794 509939 344414 524898
rect 347514 673174 348134 707162
rect 347514 672938 347546 673174
rect 347782 672938 347866 673174
rect 348102 672938 348134 673174
rect 347514 672854 348134 672938
rect 347514 672618 347546 672854
rect 347782 672618 347866 672854
rect 348102 672618 348134 672854
rect 347514 637174 348134 672618
rect 347514 636938 347546 637174
rect 347782 636938 347866 637174
rect 348102 636938 348134 637174
rect 347514 636854 348134 636938
rect 347514 636618 347546 636854
rect 347782 636618 347866 636854
rect 348102 636618 348134 636854
rect 347514 601174 348134 636618
rect 347514 600938 347546 601174
rect 347782 600938 347866 601174
rect 348102 600938 348134 601174
rect 347514 600854 348134 600938
rect 347514 600618 347546 600854
rect 347782 600618 347866 600854
rect 348102 600618 348134 600854
rect 347514 565174 348134 600618
rect 347514 564938 347546 565174
rect 347782 564938 347866 565174
rect 348102 564938 348134 565174
rect 347514 564854 348134 564938
rect 347514 564618 347546 564854
rect 347782 564618 347866 564854
rect 348102 564618 348134 564854
rect 347514 529174 348134 564618
rect 347514 528938 347546 529174
rect 347782 528938 347866 529174
rect 348102 528938 348134 529174
rect 347514 528854 348134 528938
rect 347514 528618 347546 528854
rect 347782 528618 347866 528854
rect 348102 528618 348134 528854
rect 347514 509939 348134 528618
rect 351234 676894 351854 709082
rect 351234 676658 351266 676894
rect 351502 676658 351586 676894
rect 351822 676658 351854 676894
rect 351234 676574 351854 676658
rect 351234 676338 351266 676574
rect 351502 676338 351586 676574
rect 351822 676338 351854 676574
rect 351234 640894 351854 676338
rect 351234 640658 351266 640894
rect 351502 640658 351586 640894
rect 351822 640658 351854 640894
rect 351234 640574 351854 640658
rect 351234 640338 351266 640574
rect 351502 640338 351586 640574
rect 351822 640338 351854 640574
rect 351234 604894 351854 640338
rect 351234 604658 351266 604894
rect 351502 604658 351586 604894
rect 351822 604658 351854 604894
rect 351234 604574 351854 604658
rect 351234 604338 351266 604574
rect 351502 604338 351586 604574
rect 351822 604338 351854 604574
rect 351234 568894 351854 604338
rect 351234 568658 351266 568894
rect 351502 568658 351586 568894
rect 351822 568658 351854 568894
rect 351234 568574 351854 568658
rect 351234 568338 351266 568574
rect 351502 568338 351586 568574
rect 351822 568338 351854 568574
rect 351234 532894 351854 568338
rect 351234 532658 351266 532894
rect 351502 532658 351586 532894
rect 351822 532658 351854 532894
rect 351234 532574 351854 532658
rect 351234 532338 351266 532574
rect 351502 532338 351586 532574
rect 351822 532338 351854 532574
rect 351234 509939 351854 532338
rect 354954 680614 355574 711002
rect 372954 710598 373574 711590
rect 372954 710362 372986 710598
rect 373222 710362 373306 710598
rect 373542 710362 373574 710598
rect 372954 710278 373574 710362
rect 372954 710042 372986 710278
rect 373222 710042 373306 710278
rect 373542 710042 373574 710278
rect 369234 708678 369854 709670
rect 369234 708442 369266 708678
rect 369502 708442 369586 708678
rect 369822 708442 369854 708678
rect 369234 708358 369854 708442
rect 369234 708122 369266 708358
rect 369502 708122 369586 708358
rect 369822 708122 369854 708358
rect 365514 706758 366134 707750
rect 365514 706522 365546 706758
rect 365782 706522 365866 706758
rect 366102 706522 366134 706758
rect 365514 706438 366134 706522
rect 365514 706202 365546 706438
rect 365782 706202 365866 706438
rect 366102 706202 366134 706438
rect 354954 680378 354986 680614
rect 355222 680378 355306 680614
rect 355542 680378 355574 680614
rect 354954 680294 355574 680378
rect 354954 680058 354986 680294
rect 355222 680058 355306 680294
rect 355542 680058 355574 680294
rect 354954 644614 355574 680058
rect 354954 644378 354986 644614
rect 355222 644378 355306 644614
rect 355542 644378 355574 644614
rect 354954 644294 355574 644378
rect 354954 644058 354986 644294
rect 355222 644058 355306 644294
rect 355542 644058 355574 644294
rect 354954 608614 355574 644058
rect 354954 608378 354986 608614
rect 355222 608378 355306 608614
rect 355542 608378 355574 608614
rect 354954 608294 355574 608378
rect 354954 608058 354986 608294
rect 355222 608058 355306 608294
rect 355542 608058 355574 608294
rect 354954 572614 355574 608058
rect 354954 572378 354986 572614
rect 355222 572378 355306 572614
rect 355542 572378 355574 572614
rect 354954 572294 355574 572378
rect 354954 572058 354986 572294
rect 355222 572058 355306 572294
rect 355542 572058 355574 572294
rect 354954 536614 355574 572058
rect 354954 536378 354986 536614
rect 355222 536378 355306 536614
rect 355542 536378 355574 536614
rect 354954 536294 355574 536378
rect 354954 536058 354986 536294
rect 355222 536058 355306 536294
rect 355542 536058 355574 536294
rect 354954 509939 355574 536058
rect 361794 704838 362414 705830
rect 361794 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 362414 704838
rect 361794 704518 362414 704602
rect 361794 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 362414 704518
rect 361794 687454 362414 704282
rect 361794 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 362414 687454
rect 361794 687134 362414 687218
rect 361794 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 362414 687134
rect 361794 651454 362414 686898
rect 361794 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 362414 651454
rect 361794 651134 362414 651218
rect 361794 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 362414 651134
rect 361794 615454 362414 650898
rect 361794 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 362414 615454
rect 361794 615134 362414 615218
rect 361794 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 362414 615134
rect 361794 579454 362414 614898
rect 361794 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 362414 579454
rect 361794 579134 362414 579218
rect 361794 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 362414 579134
rect 361794 543454 362414 578898
rect 361794 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 362414 543454
rect 361794 543134 362414 543218
rect 361794 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 362414 543134
rect 361794 509939 362414 542898
rect 365514 691174 366134 706202
rect 365514 690938 365546 691174
rect 365782 690938 365866 691174
rect 366102 690938 366134 691174
rect 365514 690854 366134 690938
rect 365514 690618 365546 690854
rect 365782 690618 365866 690854
rect 366102 690618 366134 690854
rect 365514 655174 366134 690618
rect 365514 654938 365546 655174
rect 365782 654938 365866 655174
rect 366102 654938 366134 655174
rect 365514 654854 366134 654938
rect 365514 654618 365546 654854
rect 365782 654618 365866 654854
rect 366102 654618 366134 654854
rect 365514 619174 366134 654618
rect 365514 618938 365546 619174
rect 365782 618938 365866 619174
rect 366102 618938 366134 619174
rect 365514 618854 366134 618938
rect 365514 618618 365546 618854
rect 365782 618618 365866 618854
rect 366102 618618 366134 618854
rect 365514 583174 366134 618618
rect 365514 582938 365546 583174
rect 365782 582938 365866 583174
rect 366102 582938 366134 583174
rect 365514 582854 366134 582938
rect 365514 582618 365546 582854
rect 365782 582618 365866 582854
rect 366102 582618 366134 582854
rect 365514 547174 366134 582618
rect 365514 546938 365546 547174
rect 365782 546938 365866 547174
rect 366102 546938 366134 547174
rect 365514 546854 366134 546938
rect 365514 546618 365546 546854
rect 365782 546618 365866 546854
rect 366102 546618 366134 546854
rect 365514 511174 366134 546618
rect 365514 510938 365546 511174
rect 365782 510938 365866 511174
rect 366102 510938 366134 511174
rect 365514 510854 366134 510938
rect 365514 510618 365546 510854
rect 365782 510618 365866 510854
rect 366102 510618 366134 510854
rect 365514 509939 366134 510618
rect 369234 694894 369854 708122
rect 369234 694658 369266 694894
rect 369502 694658 369586 694894
rect 369822 694658 369854 694894
rect 369234 694574 369854 694658
rect 369234 694338 369266 694574
rect 369502 694338 369586 694574
rect 369822 694338 369854 694574
rect 369234 658894 369854 694338
rect 369234 658658 369266 658894
rect 369502 658658 369586 658894
rect 369822 658658 369854 658894
rect 369234 658574 369854 658658
rect 369234 658338 369266 658574
rect 369502 658338 369586 658574
rect 369822 658338 369854 658574
rect 369234 622894 369854 658338
rect 369234 622658 369266 622894
rect 369502 622658 369586 622894
rect 369822 622658 369854 622894
rect 369234 622574 369854 622658
rect 369234 622338 369266 622574
rect 369502 622338 369586 622574
rect 369822 622338 369854 622574
rect 369234 586894 369854 622338
rect 369234 586658 369266 586894
rect 369502 586658 369586 586894
rect 369822 586658 369854 586894
rect 369234 586574 369854 586658
rect 369234 586338 369266 586574
rect 369502 586338 369586 586574
rect 369822 586338 369854 586574
rect 369234 550894 369854 586338
rect 369234 550658 369266 550894
rect 369502 550658 369586 550894
rect 369822 550658 369854 550894
rect 369234 550574 369854 550658
rect 369234 550338 369266 550574
rect 369502 550338 369586 550574
rect 369822 550338 369854 550574
rect 369234 514894 369854 550338
rect 369234 514658 369266 514894
rect 369502 514658 369586 514894
rect 369822 514658 369854 514894
rect 369234 514574 369854 514658
rect 369234 514338 369266 514574
rect 369502 514338 369586 514574
rect 369822 514338 369854 514574
rect 369234 509939 369854 514338
rect 372954 698614 373574 710042
rect 390954 711558 391574 711590
rect 390954 711322 390986 711558
rect 391222 711322 391306 711558
rect 391542 711322 391574 711558
rect 390954 711238 391574 711322
rect 390954 711002 390986 711238
rect 391222 711002 391306 711238
rect 391542 711002 391574 711238
rect 387234 709638 387854 709670
rect 387234 709402 387266 709638
rect 387502 709402 387586 709638
rect 387822 709402 387854 709638
rect 387234 709318 387854 709402
rect 387234 709082 387266 709318
rect 387502 709082 387586 709318
rect 387822 709082 387854 709318
rect 383514 707718 384134 707750
rect 383514 707482 383546 707718
rect 383782 707482 383866 707718
rect 384102 707482 384134 707718
rect 383514 707398 384134 707482
rect 383514 707162 383546 707398
rect 383782 707162 383866 707398
rect 384102 707162 384134 707398
rect 372954 698378 372986 698614
rect 373222 698378 373306 698614
rect 373542 698378 373574 698614
rect 372954 698294 373574 698378
rect 372954 698058 372986 698294
rect 373222 698058 373306 698294
rect 373542 698058 373574 698294
rect 372954 662614 373574 698058
rect 372954 662378 372986 662614
rect 373222 662378 373306 662614
rect 373542 662378 373574 662614
rect 372954 662294 373574 662378
rect 372954 662058 372986 662294
rect 373222 662058 373306 662294
rect 373542 662058 373574 662294
rect 372954 626614 373574 662058
rect 372954 626378 372986 626614
rect 373222 626378 373306 626614
rect 373542 626378 373574 626614
rect 372954 626294 373574 626378
rect 372954 626058 372986 626294
rect 373222 626058 373306 626294
rect 373542 626058 373574 626294
rect 372954 590614 373574 626058
rect 372954 590378 372986 590614
rect 373222 590378 373306 590614
rect 373542 590378 373574 590614
rect 372954 590294 373574 590378
rect 372954 590058 372986 590294
rect 373222 590058 373306 590294
rect 373542 590058 373574 590294
rect 372954 554614 373574 590058
rect 372954 554378 372986 554614
rect 373222 554378 373306 554614
rect 373542 554378 373574 554614
rect 372954 554294 373574 554378
rect 372954 554058 372986 554294
rect 373222 554058 373306 554294
rect 373542 554058 373574 554294
rect 372954 518614 373574 554058
rect 372954 518378 372986 518614
rect 373222 518378 373306 518614
rect 373542 518378 373574 518614
rect 372954 518294 373574 518378
rect 372954 518058 372986 518294
rect 373222 518058 373306 518294
rect 373542 518058 373574 518294
rect 372954 509939 373574 518058
rect 379794 705798 380414 705830
rect 379794 705562 379826 705798
rect 380062 705562 380146 705798
rect 380382 705562 380414 705798
rect 379794 705478 380414 705562
rect 379794 705242 379826 705478
rect 380062 705242 380146 705478
rect 380382 705242 380414 705478
rect 379794 669454 380414 705242
rect 379794 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 380414 669454
rect 379794 669134 380414 669218
rect 379794 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 380414 669134
rect 379794 633454 380414 668898
rect 379794 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 380414 633454
rect 379794 633134 380414 633218
rect 379794 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 380414 633134
rect 379794 597454 380414 632898
rect 379794 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 380414 597454
rect 379794 597134 380414 597218
rect 379794 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 380414 597134
rect 379794 561454 380414 596898
rect 379794 561218 379826 561454
rect 380062 561218 380146 561454
rect 380382 561218 380414 561454
rect 379794 561134 380414 561218
rect 379794 560898 379826 561134
rect 380062 560898 380146 561134
rect 380382 560898 380414 561134
rect 379794 525454 380414 560898
rect 379794 525218 379826 525454
rect 380062 525218 380146 525454
rect 380382 525218 380414 525454
rect 379794 525134 380414 525218
rect 379794 524898 379826 525134
rect 380062 524898 380146 525134
rect 380382 524898 380414 525134
rect 379794 509939 380414 524898
rect 383514 673174 384134 707162
rect 383514 672938 383546 673174
rect 383782 672938 383866 673174
rect 384102 672938 384134 673174
rect 383514 672854 384134 672938
rect 383514 672618 383546 672854
rect 383782 672618 383866 672854
rect 384102 672618 384134 672854
rect 383514 637174 384134 672618
rect 383514 636938 383546 637174
rect 383782 636938 383866 637174
rect 384102 636938 384134 637174
rect 383514 636854 384134 636938
rect 383514 636618 383546 636854
rect 383782 636618 383866 636854
rect 384102 636618 384134 636854
rect 383514 601174 384134 636618
rect 383514 600938 383546 601174
rect 383782 600938 383866 601174
rect 384102 600938 384134 601174
rect 383514 600854 384134 600938
rect 383514 600618 383546 600854
rect 383782 600618 383866 600854
rect 384102 600618 384134 600854
rect 383514 565174 384134 600618
rect 383514 564938 383546 565174
rect 383782 564938 383866 565174
rect 384102 564938 384134 565174
rect 383514 564854 384134 564938
rect 383514 564618 383546 564854
rect 383782 564618 383866 564854
rect 384102 564618 384134 564854
rect 383514 529174 384134 564618
rect 383514 528938 383546 529174
rect 383782 528938 383866 529174
rect 384102 528938 384134 529174
rect 383514 528854 384134 528938
rect 383514 528618 383546 528854
rect 383782 528618 383866 528854
rect 384102 528618 384134 528854
rect 383514 509939 384134 528618
rect 387234 676894 387854 709082
rect 387234 676658 387266 676894
rect 387502 676658 387586 676894
rect 387822 676658 387854 676894
rect 387234 676574 387854 676658
rect 387234 676338 387266 676574
rect 387502 676338 387586 676574
rect 387822 676338 387854 676574
rect 387234 640894 387854 676338
rect 387234 640658 387266 640894
rect 387502 640658 387586 640894
rect 387822 640658 387854 640894
rect 387234 640574 387854 640658
rect 387234 640338 387266 640574
rect 387502 640338 387586 640574
rect 387822 640338 387854 640574
rect 387234 604894 387854 640338
rect 387234 604658 387266 604894
rect 387502 604658 387586 604894
rect 387822 604658 387854 604894
rect 387234 604574 387854 604658
rect 387234 604338 387266 604574
rect 387502 604338 387586 604574
rect 387822 604338 387854 604574
rect 387234 568894 387854 604338
rect 387234 568658 387266 568894
rect 387502 568658 387586 568894
rect 387822 568658 387854 568894
rect 387234 568574 387854 568658
rect 387234 568338 387266 568574
rect 387502 568338 387586 568574
rect 387822 568338 387854 568574
rect 387234 532894 387854 568338
rect 387234 532658 387266 532894
rect 387502 532658 387586 532894
rect 387822 532658 387854 532894
rect 387234 532574 387854 532658
rect 387234 532338 387266 532574
rect 387502 532338 387586 532574
rect 387822 532338 387854 532574
rect 387234 509939 387854 532338
rect 390954 680614 391574 711002
rect 408954 710598 409574 711590
rect 408954 710362 408986 710598
rect 409222 710362 409306 710598
rect 409542 710362 409574 710598
rect 408954 710278 409574 710362
rect 408954 710042 408986 710278
rect 409222 710042 409306 710278
rect 409542 710042 409574 710278
rect 405234 708678 405854 709670
rect 405234 708442 405266 708678
rect 405502 708442 405586 708678
rect 405822 708442 405854 708678
rect 405234 708358 405854 708442
rect 405234 708122 405266 708358
rect 405502 708122 405586 708358
rect 405822 708122 405854 708358
rect 401514 706758 402134 707750
rect 401514 706522 401546 706758
rect 401782 706522 401866 706758
rect 402102 706522 402134 706758
rect 401514 706438 402134 706522
rect 401514 706202 401546 706438
rect 401782 706202 401866 706438
rect 402102 706202 402134 706438
rect 390954 680378 390986 680614
rect 391222 680378 391306 680614
rect 391542 680378 391574 680614
rect 390954 680294 391574 680378
rect 390954 680058 390986 680294
rect 391222 680058 391306 680294
rect 391542 680058 391574 680294
rect 390954 644614 391574 680058
rect 390954 644378 390986 644614
rect 391222 644378 391306 644614
rect 391542 644378 391574 644614
rect 390954 644294 391574 644378
rect 390954 644058 390986 644294
rect 391222 644058 391306 644294
rect 391542 644058 391574 644294
rect 390954 608614 391574 644058
rect 390954 608378 390986 608614
rect 391222 608378 391306 608614
rect 391542 608378 391574 608614
rect 390954 608294 391574 608378
rect 390954 608058 390986 608294
rect 391222 608058 391306 608294
rect 391542 608058 391574 608294
rect 390954 572614 391574 608058
rect 390954 572378 390986 572614
rect 391222 572378 391306 572614
rect 391542 572378 391574 572614
rect 390954 572294 391574 572378
rect 390954 572058 390986 572294
rect 391222 572058 391306 572294
rect 391542 572058 391574 572294
rect 390954 536614 391574 572058
rect 390954 536378 390986 536614
rect 391222 536378 391306 536614
rect 391542 536378 391574 536614
rect 390954 536294 391574 536378
rect 390954 536058 390986 536294
rect 391222 536058 391306 536294
rect 391542 536058 391574 536294
rect 390954 509939 391574 536058
rect 397794 704838 398414 705830
rect 397794 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 398414 704838
rect 397794 704518 398414 704602
rect 397794 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 398414 704518
rect 397794 687454 398414 704282
rect 397794 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 398414 687454
rect 397794 687134 398414 687218
rect 397794 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 398414 687134
rect 397794 651454 398414 686898
rect 397794 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 398414 651454
rect 397794 651134 398414 651218
rect 397794 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 398414 651134
rect 397794 615454 398414 650898
rect 397794 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 398414 615454
rect 397794 615134 398414 615218
rect 397794 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 398414 615134
rect 397794 579454 398414 614898
rect 397794 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 398414 579454
rect 397794 579134 398414 579218
rect 397794 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 398414 579134
rect 397794 543454 398414 578898
rect 397794 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 398414 543454
rect 397794 543134 398414 543218
rect 397794 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 398414 543134
rect 397794 509939 398414 542898
rect 401514 691174 402134 706202
rect 401514 690938 401546 691174
rect 401782 690938 401866 691174
rect 402102 690938 402134 691174
rect 401514 690854 402134 690938
rect 401514 690618 401546 690854
rect 401782 690618 401866 690854
rect 402102 690618 402134 690854
rect 401514 655174 402134 690618
rect 401514 654938 401546 655174
rect 401782 654938 401866 655174
rect 402102 654938 402134 655174
rect 401514 654854 402134 654938
rect 401514 654618 401546 654854
rect 401782 654618 401866 654854
rect 402102 654618 402134 654854
rect 401514 619174 402134 654618
rect 401514 618938 401546 619174
rect 401782 618938 401866 619174
rect 402102 618938 402134 619174
rect 401514 618854 402134 618938
rect 401514 618618 401546 618854
rect 401782 618618 401866 618854
rect 402102 618618 402134 618854
rect 401514 583174 402134 618618
rect 401514 582938 401546 583174
rect 401782 582938 401866 583174
rect 402102 582938 402134 583174
rect 401514 582854 402134 582938
rect 401514 582618 401546 582854
rect 401782 582618 401866 582854
rect 402102 582618 402134 582854
rect 401514 547174 402134 582618
rect 401514 546938 401546 547174
rect 401782 546938 401866 547174
rect 402102 546938 402134 547174
rect 401514 546854 402134 546938
rect 401514 546618 401546 546854
rect 401782 546618 401866 546854
rect 402102 546618 402134 546854
rect 401514 511174 402134 546618
rect 401514 510938 401546 511174
rect 401782 510938 401866 511174
rect 402102 510938 402134 511174
rect 401514 510854 402134 510938
rect 401514 510618 401546 510854
rect 401782 510618 401866 510854
rect 402102 510618 402134 510854
rect 401514 509939 402134 510618
rect 405234 694894 405854 708122
rect 405234 694658 405266 694894
rect 405502 694658 405586 694894
rect 405822 694658 405854 694894
rect 405234 694574 405854 694658
rect 405234 694338 405266 694574
rect 405502 694338 405586 694574
rect 405822 694338 405854 694574
rect 405234 658894 405854 694338
rect 405234 658658 405266 658894
rect 405502 658658 405586 658894
rect 405822 658658 405854 658894
rect 405234 658574 405854 658658
rect 405234 658338 405266 658574
rect 405502 658338 405586 658574
rect 405822 658338 405854 658574
rect 405234 622894 405854 658338
rect 405234 622658 405266 622894
rect 405502 622658 405586 622894
rect 405822 622658 405854 622894
rect 405234 622574 405854 622658
rect 405234 622338 405266 622574
rect 405502 622338 405586 622574
rect 405822 622338 405854 622574
rect 405234 586894 405854 622338
rect 405234 586658 405266 586894
rect 405502 586658 405586 586894
rect 405822 586658 405854 586894
rect 405234 586574 405854 586658
rect 405234 586338 405266 586574
rect 405502 586338 405586 586574
rect 405822 586338 405854 586574
rect 405234 550894 405854 586338
rect 405234 550658 405266 550894
rect 405502 550658 405586 550894
rect 405822 550658 405854 550894
rect 405234 550574 405854 550658
rect 405234 550338 405266 550574
rect 405502 550338 405586 550574
rect 405822 550338 405854 550574
rect 405234 514894 405854 550338
rect 405234 514658 405266 514894
rect 405502 514658 405586 514894
rect 405822 514658 405854 514894
rect 405234 514574 405854 514658
rect 405234 514338 405266 514574
rect 405502 514338 405586 514574
rect 405822 514338 405854 514574
rect 405234 509939 405854 514338
rect 408954 698614 409574 710042
rect 426954 711558 427574 711590
rect 426954 711322 426986 711558
rect 427222 711322 427306 711558
rect 427542 711322 427574 711558
rect 426954 711238 427574 711322
rect 426954 711002 426986 711238
rect 427222 711002 427306 711238
rect 427542 711002 427574 711238
rect 423234 709638 423854 709670
rect 423234 709402 423266 709638
rect 423502 709402 423586 709638
rect 423822 709402 423854 709638
rect 423234 709318 423854 709402
rect 423234 709082 423266 709318
rect 423502 709082 423586 709318
rect 423822 709082 423854 709318
rect 419514 707718 420134 707750
rect 419514 707482 419546 707718
rect 419782 707482 419866 707718
rect 420102 707482 420134 707718
rect 419514 707398 420134 707482
rect 419514 707162 419546 707398
rect 419782 707162 419866 707398
rect 420102 707162 420134 707398
rect 408954 698378 408986 698614
rect 409222 698378 409306 698614
rect 409542 698378 409574 698614
rect 408954 698294 409574 698378
rect 408954 698058 408986 698294
rect 409222 698058 409306 698294
rect 409542 698058 409574 698294
rect 408954 662614 409574 698058
rect 408954 662378 408986 662614
rect 409222 662378 409306 662614
rect 409542 662378 409574 662614
rect 408954 662294 409574 662378
rect 408954 662058 408986 662294
rect 409222 662058 409306 662294
rect 409542 662058 409574 662294
rect 408954 626614 409574 662058
rect 408954 626378 408986 626614
rect 409222 626378 409306 626614
rect 409542 626378 409574 626614
rect 408954 626294 409574 626378
rect 408954 626058 408986 626294
rect 409222 626058 409306 626294
rect 409542 626058 409574 626294
rect 408954 590614 409574 626058
rect 408954 590378 408986 590614
rect 409222 590378 409306 590614
rect 409542 590378 409574 590614
rect 408954 590294 409574 590378
rect 408954 590058 408986 590294
rect 409222 590058 409306 590294
rect 409542 590058 409574 590294
rect 408954 554614 409574 590058
rect 408954 554378 408986 554614
rect 409222 554378 409306 554614
rect 409542 554378 409574 554614
rect 408954 554294 409574 554378
rect 408954 554058 408986 554294
rect 409222 554058 409306 554294
rect 409542 554058 409574 554294
rect 408954 518614 409574 554058
rect 408954 518378 408986 518614
rect 409222 518378 409306 518614
rect 409542 518378 409574 518614
rect 408954 518294 409574 518378
rect 408954 518058 408986 518294
rect 409222 518058 409306 518294
rect 409542 518058 409574 518294
rect 408954 509939 409574 518058
rect 415794 705798 416414 705830
rect 415794 705562 415826 705798
rect 416062 705562 416146 705798
rect 416382 705562 416414 705798
rect 415794 705478 416414 705562
rect 415794 705242 415826 705478
rect 416062 705242 416146 705478
rect 416382 705242 416414 705478
rect 415794 669454 416414 705242
rect 415794 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 416414 669454
rect 415794 669134 416414 669218
rect 415794 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 416414 669134
rect 415794 633454 416414 668898
rect 415794 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 416414 633454
rect 415794 633134 416414 633218
rect 415794 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 416414 633134
rect 415794 597454 416414 632898
rect 415794 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 416414 597454
rect 415794 597134 416414 597218
rect 415794 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 416414 597134
rect 415794 561454 416414 596898
rect 415794 561218 415826 561454
rect 416062 561218 416146 561454
rect 416382 561218 416414 561454
rect 415794 561134 416414 561218
rect 415794 560898 415826 561134
rect 416062 560898 416146 561134
rect 416382 560898 416414 561134
rect 415794 525454 416414 560898
rect 415794 525218 415826 525454
rect 416062 525218 416146 525454
rect 416382 525218 416414 525454
rect 415794 525134 416414 525218
rect 415794 524898 415826 525134
rect 416062 524898 416146 525134
rect 416382 524898 416414 525134
rect 415794 509939 416414 524898
rect 419514 673174 420134 707162
rect 419514 672938 419546 673174
rect 419782 672938 419866 673174
rect 420102 672938 420134 673174
rect 419514 672854 420134 672938
rect 419514 672618 419546 672854
rect 419782 672618 419866 672854
rect 420102 672618 420134 672854
rect 419514 637174 420134 672618
rect 419514 636938 419546 637174
rect 419782 636938 419866 637174
rect 420102 636938 420134 637174
rect 419514 636854 420134 636938
rect 419514 636618 419546 636854
rect 419782 636618 419866 636854
rect 420102 636618 420134 636854
rect 419514 601174 420134 636618
rect 419514 600938 419546 601174
rect 419782 600938 419866 601174
rect 420102 600938 420134 601174
rect 419514 600854 420134 600938
rect 419514 600618 419546 600854
rect 419782 600618 419866 600854
rect 420102 600618 420134 600854
rect 419514 565174 420134 600618
rect 419514 564938 419546 565174
rect 419782 564938 419866 565174
rect 420102 564938 420134 565174
rect 419514 564854 420134 564938
rect 419514 564618 419546 564854
rect 419782 564618 419866 564854
rect 420102 564618 420134 564854
rect 419514 529174 420134 564618
rect 419514 528938 419546 529174
rect 419782 528938 419866 529174
rect 420102 528938 420134 529174
rect 419514 528854 420134 528938
rect 419514 528618 419546 528854
rect 419782 528618 419866 528854
rect 420102 528618 420134 528854
rect 419514 509939 420134 528618
rect 423234 676894 423854 709082
rect 423234 676658 423266 676894
rect 423502 676658 423586 676894
rect 423822 676658 423854 676894
rect 423234 676574 423854 676658
rect 423234 676338 423266 676574
rect 423502 676338 423586 676574
rect 423822 676338 423854 676574
rect 423234 640894 423854 676338
rect 423234 640658 423266 640894
rect 423502 640658 423586 640894
rect 423822 640658 423854 640894
rect 423234 640574 423854 640658
rect 423234 640338 423266 640574
rect 423502 640338 423586 640574
rect 423822 640338 423854 640574
rect 423234 604894 423854 640338
rect 423234 604658 423266 604894
rect 423502 604658 423586 604894
rect 423822 604658 423854 604894
rect 423234 604574 423854 604658
rect 423234 604338 423266 604574
rect 423502 604338 423586 604574
rect 423822 604338 423854 604574
rect 423234 568894 423854 604338
rect 423234 568658 423266 568894
rect 423502 568658 423586 568894
rect 423822 568658 423854 568894
rect 423234 568574 423854 568658
rect 423234 568338 423266 568574
rect 423502 568338 423586 568574
rect 423822 568338 423854 568574
rect 423234 532894 423854 568338
rect 423234 532658 423266 532894
rect 423502 532658 423586 532894
rect 423822 532658 423854 532894
rect 423234 532574 423854 532658
rect 423234 532338 423266 532574
rect 423502 532338 423586 532574
rect 423822 532338 423854 532574
rect 423234 496894 423854 532338
rect 423234 496658 423266 496894
rect 423502 496658 423586 496894
rect 423822 496658 423854 496894
rect 423234 496574 423854 496658
rect 423234 496338 423266 496574
rect 423502 496338 423586 496574
rect 423822 496338 423854 496574
rect 185368 489454 185688 489486
rect 185368 489218 185410 489454
rect 185646 489218 185688 489454
rect 185368 489134 185688 489218
rect 185368 488898 185410 489134
rect 185646 488898 185688 489134
rect 185368 488866 185688 488898
rect 216088 489454 216408 489486
rect 216088 489218 216130 489454
rect 216366 489218 216408 489454
rect 216088 489134 216408 489218
rect 216088 488898 216130 489134
rect 216366 488898 216408 489134
rect 216088 488866 216408 488898
rect 246808 489454 247128 489486
rect 246808 489218 246850 489454
rect 247086 489218 247128 489454
rect 246808 489134 247128 489218
rect 246808 488898 246850 489134
rect 247086 488898 247128 489134
rect 246808 488866 247128 488898
rect 277528 489454 277848 489486
rect 277528 489218 277570 489454
rect 277806 489218 277848 489454
rect 277528 489134 277848 489218
rect 277528 488898 277570 489134
rect 277806 488898 277848 489134
rect 277528 488866 277848 488898
rect 308248 489454 308568 489486
rect 308248 489218 308290 489454
rect 308526 489218 308568 489454
rect 308248 489134 308568 489218
rect 308248 488898 308290 489134
rect 308526 488898 308568 489134
rect 308248 488866 308568 488898
rect 338968 489454 339288 489486
rect 338968 489218 339010 489454
rect 339246 489218 339288 489454
rect 338968 489134 339288 489218
rect 338968 488898 339010 489134
rect 339246 488898 339288 489134
rect 338968 488866 339288 488898
rect 369688 489454 370008 489486
rect 369688 489218 369730 489454
rect 369966 489218 370008 489454
rect 369688 489134 370008 489218
rect 369688 488898 369730 489134
rect 369966 488898 370008 489134
rect 369688 488866 370008 488898
rect 400408 489454 400728 489486
rect 400408 489218 400450 489454
rect 400686 489218 400728 489454
rect 400408 489134 400728 489218
rect 400408 488898 400450 489134
rect 400686 488898 400728 489134
rect 400408 488866 400728 488898
rect 156954 482378 156986 482614
rect 157222 482378 157306 482614
rect 157542 482378 157574 482614
rect 156954 482294 157574 482378
rect 156954 482058 156986 482294
rect 157222 482058 157306 482294
rect 157542 482058 157574 482294
rect 156954 446614 157574 482058
rect 170008 471454 170328 471486
rect 170008 471218 170050 471454
rect 170286 471218 170328 471454
rect 170008 471134 170328 471218
rect 170008 470898 170050 471134
rect 170286 470898 170328 471134
rect 170008 470866 170328 470898
rect 200728 471454 201048 471486
rect 200728 471218 200770 471454
rect 201006 471218 201048 471454
rect 200728 471134 201048 471218
rect 200728 470898 200770 471134
rect 201006 470898 201048 471134
rect 200728 470866 201048 470898
rect 231448 471454 231768 471486
rect 231448 471218 231490 471454
rect 231726 471218 231768 471454
rect 231448 471134 231768 471218
rect 231448 470898 231490 471134
rect 231726 470898 231768 471134
rect 231448 470866 231768 470898
rect 262168 471454 262488 471486
rect 262168 471218 262210 471454
rect 262446 471218 262488 471454
rect 262168 471134 262488 471218
rect 262168 470898 262210 471134
rect 262446 470898 262488 471134
rect 262168 470866 262488 470898
rect 292888 471454 293208 471486
rect 292888 471218 292930 471454
rect 293166 471218 293208 471454
rect 292888 471134 293208 471218
rect 292888 470898 292930 471134
rect 293166 470898 293208 471134
rect 292888 470866 293208 470898
rect 323608 471454 323928 471486
rect 323608 471218 323650 471454
rect 323886 471218 323928 471454
rect 323608 471134 323928 471218
rect 323608 470898 323650 471134
rect 323886 470898 323928 471134
rect 323608 470866 323928 470898
rect 354328 471454 354648 471486
rect 354328 471218 354370 471454
rect 354606 471218 354648 471454
rect 354328 471134 354648 471218
rect 354328 470898 354370 471134
rect 354606 470898 354648 471134
rect 354328 470866 354648 470898
rect 385048 471454 385368 471486
rect 385048 471218 385090 471454
rect 385326 471218 385368 471454
rect 385048 471134 385368 471218
rect 385048 470898 385090 471134
rect 385326 470898 385368 471134
rect 385048 470866 385368 470898
rect 415768 471454 416088 471486
rect 415768 471218 415810 471454
rect 416046 471218 416088 471454
rect 415768 471134 416088 471218
rect 415768 470898 415810 471134
rect 416046 470898 416088 471134
rect 415768 470866 416088 470898
rect 423234 460894 423854 496338
rect 423234 460658 423266 460894
rect 423502 460658 423586 460894
rect 423822 460658 423854 460894
rect 423234 460574 423854 460658
rect 423234 460338 423266 460574
rect 423502 460338 423586 460574
rect 423822 460338 423854 460574
rect 185368 453454 185688 453486
rect 185368 453218 185410 453454
rect 185646 453218 185688 453454
rect 185368 453134 185688 453218
rect 185368 452898 185410 453134
rect 185646 452898 185688 453134
rect 185368 452866 185688 452898
rect 216088 453454 216408 453486
rect 216088 453218 216130 453454
rect 216366 453218 216408 453454
rect 216088 453134 216408 453218
rect 216088 452898 216130 453134
rect 216366 452898 216408 453134
rect 216088 452866 216408 452898
rect 246808 453454 247128 453486
rect 246808 453218 246850 453454
rect 247086 453218 247128 453454
rect 246808 453134 247128 453218
rect 246808 452898 246850 453134
rect 247086 452898 247128 453134
rect 246808 452866 247128 452898
rect 277528 453454 277848 453486
rect 277528 453218 277570 453454
rect 277806 453218 277848 453454
rect 277528 453134 277848 453218
rect 277528 452898 277570 453134
rect 277806 452898 277848 453134
rect 277528 452866 277848 452898
rect 308248 453454 308568 453486
rect 308248 453218 308290 453454
rect 308526 453218 308568 453454
rect 308248 453134 308568 453218
rect 308248 452898 308290 453134
rect 308526 452898 308568 453134
rect 308248 452866 308568 452898
rect 338968 453454 339288 453486
rect 338968 453218 339010 453454
rect 339246 453218 339288 453454
rect 338968 453134 339288 453218
rect 338968 452898 339010 453134
rect 339246 452898 339288 453134
rect 338968 452866 339288 452898
rect 369688 453454 370008 453486
rect 369688 453218 369730 453454
rect 369966 453218 370008 453454
rect 369688 453134 370008 453218
rect 369688 452898 369730 453134
rect 369966 452898 370008 453134
rect 369688 452866 370008 452898
rect 400408 453454 400728 453486
rect 400408 453218 400450 453454
rect 400686 453218 400728 453454
rect 400408 453134 400728 453218
rect 400408 452898 400450 453134
rect 400686 452898 400728 453134
rect 400408 452866 400728 452898
rect 156954 446378 156986 446614
rect 157222 446378 157306 446614
rect 157542 446378 157574 446614
rect 156954 446294 157574 446378
rect 156954 446058 156986 446294
rect 157222 446058 157306 446294
rect 157542 446058 157574 446294
rect 156954 410614 157574 446058
rect 170008 435454 170328 435486
rect 170008 435218 170050 435454
rect 170286 435218 170328 435454
rect 170008 435134 170328 435218
rect 170008 434898 170050 435134
rect 170286 434898 170328 435134
rect 170008 434866 170328 434898
rect 200728 435454 201048 435486
rect 200728 435218 200770 435454
rect 201006 435218 201048 435454
rect 200728 435134 201048 435218
rect 200728 434898 200770 435134
rect 201006 434898 201048 435134
rect 200728 434866 201048 434898
rect 231448 435454 231768 435486
rect 231448 435218 231490 435454
rect 231726 435218 231768 435454
rect 231448 435134 231768 435218
rect 231448 434898 231490 435134
rect 231726 434898 231768 435134
rect 231448 434866 231768 434898
rect 262168 435454 262488 435486
rect 262168 435218 262210 435454
rect 262446 435218 262488 435454
rect 262168 435134 262488 435218
rect 262168 434898 262210 435134
rect 262446 434898 262488 435134
rect 262168 434866 262488 434898
rect 292888 435454 293208 435486
rect 292888 435218 292930 435454
rect 293166 435218 293208 435454
rect 292888 435134 293208 435218
rect 292888 434898 292930 435134
rect 293166 434898 293208 435134
rect 292888 434866 293208 434898
rect 323608 435454 323928 435486
rect 323608 435218 323650 435454
rect 323886 435218 323928 435454
rect 323608 435134 323928 435218
rect 323608 434898 323650 435134
rect 323886 434898 323928 435134
rect 323608 434866 323928 434898
rect 354328 435454 354648 435486
rect 354328 435218 354370 435454
rect 354606 435218 354648 435454
rect 354328 435134 354648 435218
rect 354328 434898 354370 435134
rect 354606 434898 354648 435134
rect 354328 434866 354648 434898
rect 385048 435454 385368 435486
rect 385048 435218 385090 435454
rect 385326 435218 385368 435454
rect 385048 435134 385368 435218
rect 385048 434898 385090 435134
rect 385326 434898 385368 435134
rect 385048 434866 385368 434898
rect 415768 435454 416088 435486
rect 415768 435218 415810 435454
rect 416046 435218 416088 435454
rect 415768 435134 416088 435218
rect 415768 434898 415810 435134
rect 416046 434898 416088 435134
rect 415768 434866 416088 434898
rect 423234 424894 423854 460338
rect 423234 424658 423266 424894
rect 423502 424658 423586 424894
rect 423822 424658 423854 424894
rect 423234 424574 423854 424658
rect 423234 424338 423266 424574
rect 423502 424338 423586 424574
rect 423822 424338 423854 424574
rect 185368 417454 185688 417486
rect 185368 417218 185410 417454
rect 185646 417218 185688 417454
rect 185368 417134 185688 417218
rect 185368 416898 185410 417134
rect 185646 416898 185688 417134
rect 185368 416866 185688 416898
rect 216088 417454 216408 417486
rect 216088 417218 216130 417454
rect 216366 417218 216408 417454
rect 216088 417134 216408 417218
rect 216088 416898 216130 417134
rect 216366 416898 216408 417134
rect 216088 416866 216408 416898
rect 246808 417454 247128 417486
rect 246808 417218 246850 417454
rect 247086 417218 247128 417454
rect 246808 417134 247128 417218
rect 246808 416898 246850 417134
rect 247086 416898 247128 417134
rect 246808 416866 247128 416898
rect 277528 417454 277848 417486
rect 277528 417218 277570 417454
rect 277806 417218 277848 417454
rect 277528 417134 277848 417218
rect 277528 416898 277570 417134
rect 277806 416898 277848 417134
rect 277528 416866 277848 416898
rect 308248 417454 308568 417486
rect 308248 417218 308290 417454
rect 308526 417218 308568 417454
rect 308248 417134 308568 417218
rect 308248 416898 308290 417134
rect 308526 416898 308568 417134
rect 308248 416866 308568 416898
rect 338968 417454 339288 417486
rect 338968 417218 339010 417454
rect 339246 417218 339288 417454
rect 338968 417134 339288 417218
rect 338968 416898 339010 417134
rect 339246 416898 339288 417134
rect 338968 416866 339288 416898
rect 369688 417454 370008 417486
rect 369688 417218 369730 417454
rect 369966 417218 370008 417454
rect 369688 417134 370008 417218
rect 369688 416898 369730 417134
rect 369966 416898 370008 417134
rect 369688 416866 370008 416898
rect 400408 417454 400728 417486
rect 400408 417218 400450 417454
rect 400686 417218 400728 417454
rect 400408 417134 400728 417218
rect 400408 416898 400450 417134
rect 400686 416898 400728 417134
rect 400408 416866 400728 416898
rect 156954 410378 156986 410614
rect 157222 410378 157306 410614
rect 157542 410378 157574 410614
rect 156954 410294 157574 410378
rect 156954 410058 156986 410294
rect 157222 410058 157306 410294
rect 157542 410058 157574 410294
rect 156954 374614 157574 410058
rect 170008 399454 170328 399486
rect 170008 399218 170050 399454
rect 170286 399218 170328 399454
rect 170008 399134 170328 399218
rect 170008 398898 170050 399134
rect 170286 398898 170328 399134
rect 170008 398866 170328 398898
rect 200728 399454 201048 399486
rect 200728 399218 200770 399454
rect 201006 399218 201048 399454
rect 200728 399134 201048 399218
rect 200728 398898 200770 399134
rect 201006 398898 201048 399134
rect 200728 398866 201048 398898
rect 231448 399454 231768 399486
rect 231448 399218 231490 399454
rect 231726 399218 231768 399454
rect 231448 399134 231768 399218
rect 231448 398898 231490 399134
rect 231726 398898 231768 399134
rect 231448 398866 231768 398898
rect 262168 399454 262488 399486
rect 262168 399218 262210 399454
rect 262446 399218 262488 399454
rect 262168 399134 262488 399218
rect 262168 398898 262210 399134
rect 262446 398898 262488 399134
rect 262168 398866 262488 398898
rect 292888 399454 293208 399486
rect 292888 399218 292930 399454
rect 293166 399218 293208 399454
rect 292888 399134 293208 399218
rect 292888 398898 292930 399134
rect 293166 398898 293208 399134
rect 292888 398866 293208 398898
rect 323608 399454 323928 399486
rect 323608 399218 323650 399454
rect 323886 399218 323928 399454
rect 323608 399134 323928 399218
rect 323608 398898 323650 399134
rect 323886 398898 323928 399134
rect 323608 398866 323928 398898
rect 354328 399454 354648 399486
rect 354328 399218 354370 399454
rect 354606 399218 354648 399454
rect 354328 399134 354648 399218
rect 354328 398898 354370 399134
rect 354606 398898 354648 399134
rect 354328 398866 354648 398898
rect 385048 399454 385368 399486
rect 385048 399218 385090 399454
rect 385326 399218 385368 399454
rect 385048 399134 385368 399218
rect 385048 398898 385090 399134
rect 385326 398898 385368 399134
rect 385048 398866 385368 398898
rect 415768 399454 416088 399486
rect 415768 399218 415810 399454
rect 416046 399218 416088 399454
rect 415768 399134 416088 399218
rect 415768 398898 415810 399134
rect 416046 398898 416088 399134
rect 415768 398866 416088 398898
rect 423234 388894 423854 424338
rect 423234 388658 423266 388894
rect 423502 388658 423586 388894
rect 423822 388658 423854 388894
rect 423234 388574 423854 388658
rect 423234 388338 423266 388574
rect 423502 388338 423586 388574
rect 423822 388338 423854 388574
rect 185368 381454 185688 381486
rect 185368 381218 185410 381454
rect 185646 381218 185688 381454
rect 185368 381134 185688 381218
rect 185368 380898 185410 381134
rect 185646 380898 185688 381134
rect 185368 380866 185688 380898
rect 216088 381454 216408 381486
rect 216088 381218 216130 381454
rect 216366 381218 216408 381454
rect 216088 381134 216408 381218
rect 216088 380898 216130 381134
rect 216366 380898 216408 381134
rect 216088 380866 216408 380898
rect 246808 381454 247128 381486
rect 246808 381218 246850 381454
rect 247086 381218 247128 381454
rect 246808 381134 247128 381218
rect 246808 380898 246850 381134
rect 247086 380898 247128 381134
rect 246808 380866 247128 380898
rect 277528 381454 277848 381486
rect 277528 381218 277570 381454
rect 277806 381218 277848 381454
rect 277528 381134 277848 381218
rect 277528 380898 277570 381134
rect 277806 380898 277848 381134
rect 277528 380866 277848 380898
rect 308248 381454 308568 381486
rect 308248 381218 308290 381454
rect 308526 381218 308568 381454
rect 308248 381134 308568 381218
rect 308248 380898 308290 381134
rect 308526 380898 308568 381134
rect 308248 380866 308568 380898
rect 338968 381454 339288 381486
rect 338968 381218 339010 381454
rect 339246 381218 339288 381454
rect 338968 381134 339288 381218
rect 338968 380898 339010 381134
rect 339246 380898 339288 381134
rect 338968 380866 339288 380898
rect 369688 381454 370008 381486
rect 369688 381218 369730 381454
rect 369966 381218 370008 381454
rect 369688 381134 370008 381218
rect 369688 380898 369730 381134
rect 369966 380898 370008 381134
rect 369688 380866 370008 380898
rect 400408 381454 400728 381486
rect 400408 381218 400450 381454
rect 400686 381218 400728 381454
rect 400408 381134 400728 381218
rect 400408 380898 400450 381134
rect 400686 380898 400728 381134
rect 400408 380866 400728 380898
rect 156954 374378 156986 374614
rect 157222 374378 157306 374614
rect 157542 374378 157574 374614
rect 156954 374294 157574 374378
rect 156954 374058 156986 374294
rect 157222 374058 157306 374294
rect 157542 374058 157574 374294
rect 156954 338614 157574 374058
rect 170008 363454 170328 363486
rect 170008 363218 170050 363454
rect 170286 363218 170328 363454
rect 170008 363134 170328 363218
rect 170008 362898 170050 363134
rect 170286 362898 170328 363134
rect 170008 362866 170328 362898
rect 200728 363454 201048 363486
rect 200728 363218 200770 363454
rect 201006 363218 201048 363454
rect 200728 363134 201048 363218
rect 200728 362898 200770 363134
rect 201006 362898 201048 363134
rect 200728 362866 201048 362898
rect 231448 363454 231768 363486
rect 231448 363218 231490 363454
rect 231726 363218 231768 363454
rect 231448 363134 231768 363218
rect 231448 362898 231490 363134
rect 231726 362898 231768 363134
rect 231448 362866 231768 362898
rect 262168 363454 262488 363486
rect 262168 363218 262210 363454
rect 262446 363218 262488 363454
rect 262168 363134 262488 363218
rect 262168 362898 262210 363134
rect 262446 362898 262488 363134
rect 262168 362866 262488 362898
rect 292888 363454 293208 363486
rect 292888 363218 292930 363454
rect 293166 363218 293208 363454
rect 292888 363134 293208 363218
rect 292888 362898 292930 363134
rect 293166 362898 293208 363134
rect 292888 362866 293208 362898
rect 323608 363454 323928 363486
rect 323608 363218 323650 363454
rect 323886 363218 323928 363454
rect 323608 363134 323928 363218
rect 323608 362898 323650 363134
rect 323886 362898 323928 363134
rect 323608 362866 323928 362898
rect 354328 363454 354648 363486
rect 354328 363218 354370 363454
rect 354606 363218 354648 363454
rect 354328 363134 354648 363218
rect 354328 362898 354370 363134
rect 354606 362898 354648 363134
rect 354328 362866 354648 362898
rect 385048 363454 385368 363486
rect 385048 363218 385090 363454
rect 385326 363218 385368 363454
rect 385048 363134 385368 363218
rect 385048 362898 385090 363134
rect 385326 362898 385368 363134
rect 385048 362866 385368 362898
rect 415768 363454 416088 363486
rect 415768 363218 415810 363454
rect 416046 363218 416088 363454
rect 415768 363134 416088 363218
rect 415768 362898 415810 363134
rect 416046 362898 416088 363134
rect 415768 362866 416088 362898
rect 423234 352894 423854 388338
rect 423234 352658 423266 352894
rect 423502 352658 423586 352894
rect 423822 352658 423854 352894
rect 423234 352574 423854 352658
rect 423234 352338 423266 352574
rect 423502 352338 423586 352574
rect 423822 352338 423854 352574
rect 185368 345454 185688 345486
rect 185368 345218 185410 345454
rect 185646 345218 185688 345454
rect 185368 345134 185688 345218
rect 185368 344898 185410 345134
rect 185646 344898 185688 345134
rect 185368 344866 185688 344898
rect 216088 345454 216408 345486
rect 216088 345218 216130 345454
rect 216366 345218 216408 345454
rect 216088 345134 216408 345218
rect 216088 344898 216130 345134
rect 216366 344898 216408 345134
rect 216088 344866 216408 344898
rect 246808 345454 247128 345486
rect 246808 345218 246850 345454
rect 247086 345218 247128 345454
rect 246808 345134 247128 345218
rect 246808 344898 246850 345134
rect 247086 344898 247128 345134
rect 246808 344866 247128 344898
rect 277528 345454 277848 345486
rect 277528 345218 277570 345454
rect 277806 345218 277848 345454
rect 277528 345134 277848 345218
rect 277528 344898 277570 345134
rect 277806 344898 277848 345134
rect 277528 344866 277848 344898
rect 308248 345454 308568 345486
rect 308248 345218 308290 345454
rect 308526 345218 308568 345454
rect 308248 345134 308568 345218
rect 308248 344898 308290 345134
rect 308526 344898 308568 345134
rect 308248 344866 308568 344898
rect 338968 345454 339288 345486
rect 338968 345218 339010 345454
rect 339246 345218 339288 345454
rect 338968 345134 339288 345218
rect 338968 344898 339010 345134
rect 339246 344898 339288 345134
rect 338968 344866 339288 344898
rect 369688 345454 370008 345486
rect 369688 345218 369730 345454
rect 369966 345218 370008 345454
rect 369688 345134 370008 345218
rect 369688 344898 369730 345134
rect 369966 344898 370008 345134
rect 369688 344866 370008 344898
rect 400408 345454 400728 345486
rect 400408 345218 400450 345454
rect 400686 345218 400728 345454
rect 400408 345134 400728 345218
rect 400408 344898 400450 345134
rect 400686 344898 400728 345134
rect 400408 344866 400728 344898
rect 156954 338378 156986 338614
rect 157222 338378 157306 338614
rect 157542 338378 157574 338614
rect 156954 338294 157574 338378
rect 156954 338058 156986 338294
rect 157222 338058 157306 338294
rect 157542 338058 157574 338294
rect 156954 302614 157574 338058
rect 170008 327454 170328 327486
rect 170008 327218 170050 327454
rect 170286 327218 170328 327454
rect 170008 327134 170328 327218
rect 170008 326898 170050 327134
rect 170286 326898 170328 327134
rect 170008 326866 170328 326898
rect 200728 327454 201048 327486
rect 200728 327218 200770 327454
rect 201006 327218 201048 327454
rect 200728 327134 201048 327218
rect 200728 326898 200770 327134
rect 201006 326898 201048 327134
rect 200728 326866 201048 326898
rect 231448 327454 231768 327486
rect 231448 327218 231490 327454
rect 231726 327218 231768 327454
rect 231448 327134 231768 327218
rect 231448 326898 231490 327134
rect 231726 326898 231768 327134
rect 231448 326866 231768 326898
rect 262168 327454 262488 327486
rect 262168 327218 262210 327454
rect 262446 327218 262488 327454
rect 262168 327134 262488 327218
rect 262168 326898 262210 327134
rect 262446 326898 262488 327134
rect 262168 326866 262488 326898
rect 292888 327454 293208 327486
rect 292888 327218 292930 327454
rect 293166 327218 293208 327454
rect 292888 327134 293208 327218
rect 292888 326898 292930 327134
rect 293166 326898 293208 327134
rect 292888 326866 293208 326898
rect 323608 327454 323928 327486
rect 323608 327218 323650 327454
rect 323886 327218 323928 327454
rect 323608 327134 323928 327218
rect 323608 326898 323650 327134
rect 323886 326898 323928 327134
rect 323608 326866 323928 326898
rect 354328 327454 354648 327486
rect 354328 327218 354370 327454
rect 354606 327218 354648 327454
rect 354328 327134 354648 327218
rect 354328 326898 354370 327134
rect 354606 326898 354648 327134
rect 354328 326866 354648 326898
rect 385048 327454 385368 327486
rect 385048 327218 385090 327454
rect 385326 327218 385368 327454
rect 385048 327134 385368 327218
rect 385048 326898 385090 327134
rect 385326 326898 385368 327134
rect 385048 326866 385368 326898
rect 415768 327454 416088 327486
rect 415768 327218 415810 327454
rect 416046 327218 416088 327454
rect 415768 327134 416088 327218
rect 415768 326898 415810 327134
rect 416046 326898 416088 327134
rect 415768 326866 416088 326898
rect 423234 316894 423854 352338
rect 423234 316658 423266 316894
rect 423502 316658 423586 316894
rect 423822 316658 423854 316894
rect 423234 316574 423854 316658
rect 423234 316338 423266 316574
rect 423502 316338 423586 316574
rect 423822 316338 423854 316574
rect 185368 309454 185688 309486
rect 185368 309218 185410 309454
rect 185646 309218 185688 309454
rect 185368 309134 185688 309218
rect 185368 308898 185410 309134
rect 185646 308898 185688 309134
rect 185368 308866 185688 308898
rect 216088 309454 216408 309486
rect 216088 309218 216130 309454
rect 216366 309218 216408 309454
rect 216088 309134 216408 309218
rect 216088 308898 216130 309134
rect 216366 308898 216408 309134
rect 216088 308866 216408 308898
rect 246808 309454 247128 309486
rect 246808 309218 246850 309454
rect 247086 309218 247128 309454
rect 246808 309134 247128 309218
rect 246808 308898 246850 309134
rect 247086 308898 247128 309134
rect 246808 308866 247128 308898
rect 277528 309454 277848 309486
rect 277528 309218 277570 309454
rect 277806 309218 277848 309454
rect 277528 309134 277848 309218
rect 277528 308898 277570 309134
rect 277806 308898 277848 309134
rect 277528 308866 277848 308898
rect 308248 309454 308568 309486
rect 308248 309218 308290 309454
rect 308526 309218 308568 309454
rect 308248 309134 308568 309218
rect 308248 308898 308290 309134
rect 308526 308898 308568 309134
rect 308248 308866 308568 308898
rect 338968 309454 339288 309486
rect 338968 309218 339010 309454
rect 339246 309218 339288 309454
rect 338968 309134 339288 309218
rect 338968 308898 339010 309134
rect 339246 308898 339288 309134
rect 338968 308866 339288 308898
rect 369688 309454 370008 309486
rect 369688 309218 369730 309454
rect 369966 309218 370008 309454
rect 369688 309134 370008 309218
rect 369688 308898 369730 309134
rect 369966 308898 370008 309134
rect 369688 308866 370008 308898
rect 400408 309454 400728 309486
rect 400408 309218 400450 309454
rect 400686 309218 400728 309454
rect 400408 309134 400728 309218
rect 400408 308898 400450 309134
rect 400686 308898 400728 309134
rect 400408 308866 400728 308898
rect 156954 302378 156986 302614
rect 157222 302378 157306 302614
rect 157542 302378 157574 302614
rect 156954 302294 157574 302378
rect 156954 302058 156986 302294
rect 157222 302058 157306 302294
rect 157542 302058 157574 302294
rect 156954 266614 157574 302058
rect 170008 291454 170328 291486
rect 170008 291218 170050 291454
rect 170286 291218 170328 291454
rect 170008 291134 170328 291218
rect 170008 290898 170050 291134
rect 170286 290898 170328 291134
rect 170008 290866 170328 290898
rect 200728 291454 201048 291486
rect 200728 291218 200770 291454
rect 201006 291218 201048 291454
rect 200728 291134 201048 291218
rect 200728 290898 200770 291134
rect 201006 290898 201048 291134
rect 200728 290866 201048 290898
rect 231448 291454 231768 291486
rect 231448 291218 231490 291454
rect 231726 291218 231768 291454
rect 231448 291134 231768 291218
rect 231448 290898 231490 291134
rect 231726 290898 231768 291134
rect 231448 290866 231768 290898
rect 262168 291454 262488 291486
rect 262168 291218 262210 291454
rect 262446 291218 262488 291454
rect 262168 291134 262488 291218
rect 262168 290898 262210 291134
rect 262446 290898 262488 291134
rect 262168 290866 262488 290898
rect 292888 291454 293208 291486
rect 292888 291218 292930 291454
rect 293166 291218 293208 291454
rect 292888 291134 293208 291218
rect 292888 290898 292930 291134
rect 293166 290898 293208 291134
rect 292888 290866 293208 290898
rect 323608 291454 323928 291486
rect 323608 291218 323650 291454
rect 323886 291218 323928 291454
rect 323608 291134 323928 291218
rect 323608 290898 323650 291134
rect 323886 290898 323928 291134
rect 323608 290866 323928 290898
rect 354328 291454 354648 291486
rect 354328 291218 354370 291454
rect 354606 291218 354648 291454
rect 354328 291134 354648 291218
rect 354328 290898 354370 291134
rect 354606 290898 354648 291134
rect 354328 290866 354648 290898
rect 385048 291454 385368 291486
rect 385048 291218 385090 291454
rect 385326 291218 385368 291454
rect 385048 291134 385368 291218
rect 385048 290898 385090 291134
rect 385326 290898 385368 291134
rect 385048 290866 385368 290898
rect 415768 291454 416088 291486
rect 415768 291218 415810 291454
rect 416046 291218 416088 291454
rect 415768 291134 416088 291218
rect 415768 290898 415810 291134
rect 416046 290898 416088 291134
rect 415768 290866 416088 290898
rect 423234 280894 423854 316338
rect 423234 280658 423266 280894
rect 423502 280658 423586 280894
rect 423822 280658 423854 280894
rect 423234 280574 423854 280658
rect 423234 280338 423266 280574
rect 423502 280338 423586 280574
rect 423822 280338 423854 280574
rect 185368 273454 185688 273486
rect 185368 273218 185410 273454
rect 185646 273218 185688 273454
rect 185368 273134 185688 273218
rect 185368 272898 185410 273134
rect 185646 272898 185688 273134
rect 185368 272866 185688 272898
rect 216088 273454 216408 273486
rect 216088 273218 216130 273454
rect 216366 273218 216408 273454
rect 216088 273134 216408 273218
rect 216088 272898 216130 273134
rect 216366 272898 216408 273134
rect 216088 272866 216408 272898
rect 246808 273454 247128 273486
rect 246808 273218 246850 273454
rect 247086 273218 247128 273454
rect 246808 273134 247128 273218
rect 246808 272898 246850 273134
rect 247086 272898 247128 273134
rect 246808 272866 247128 272898
rect 277528 273454 277848 273486
rect 277528 273218 277570 273454
rect 277806 273218 277848 273454
rect 277528 273134 277848 273218
rect 277528 272898 277570 273134
rect 277806 272898 277848 273134
rect 277528 272866 277848 272898
rect 308248 273454 308568 273486
rect 308248 273218 308290 273454
rect 308526 273218 308568 273454
rect 308248 273134 308568 273218
rect 308248 272898 308290 273134
rect 308526 272898 308568 273134
rect 308248 272866 308568 272898
rect 338968 273454 339288 273486
rect 338968 273218 339010 273454
rect 339246 273218 339288 273454
rect 338968 273134 339288 273218
rect 338968 272898 339010 273134
rect 339246 272898 339288 273134
rect 338968 272866 339288 272898
rect 369688 273454 370008 273486
rect 369688 273218 369730 273454
rect 369966 273218 370008 273454
rect 369688 273134 370008 273218
rect 369688 272898 369730 273134
rect 369966 272898 370008 273134
rect 369688 272866 370008 272898
rect 400408 273454 400728 273486
rect 400408 273218 400450 273454
rect 400686 273218 400728 273454
rect 400408 273134 400728 273218
rect 400408 272898 400450 273134
rect 400686 272898 400728 273134
rect 400408 272866 400728 272898
rect 156954 266378 156986 266614
rect 157222 266378 157306 266614
rect 157542 266378 157574 266614
rect 156954 266294 157574 266378
rect 156954 266058 156986 266294
rect 157222 266058 157306 266294
rect 157542 266058 157574 266294
rect 156954 230614 157574 266058
rect 170008 255454 170328 255486
rect 170008 255218 170050 255454
rect 170286 255218 170328 255454
rect 170008 255134 170328 255218
rect 170008 254898 170050 255134
rect 170286 254898 170328 255134
rect 170008 254866 170328 254898
rect 200728 255454 201048 255486
rect 200728 255218 200770 255454
rect 201006 255218 201048 255454
rect 200728 255134 201048 255218
rect 200728 254898 200770 255134
rect 201006 254898 201048 255134
rect 200728 254866 201048 254898
rect 231448 255454 231768 255486
rect 231448 255218 231490 255454
rect 231726 255218 231768 255454
rect 231448 255134 231768 255218
rect 231448 254898 231490 255134
rect 231726 254898 231768 255134
rect 231448 254866 231768 254898
rect 262168 255454 262488 255486
rect 262168 255218 262210 255454
rect 262446 255218 262488 255454
rect 262168 255134 262488 255218
rect 262168 254898 262210 255134
rect 262446 254898 262488 255134
rect 262168 254866 262488 254898
rect 292888 255454 293208 255486
rect 292888 255218 292930 255454
rect 293166 255218 293208 255454
rect 292888 255134 293208 255218
rect 292888 254898 292930 255134
rect 293166 254898 293208 255134
rect 292888 254866 293208 254898
rect 323608 255454 323928 255486
rect 323608 255218 323650 255454
rect 323886 255218 323928 255454
rect 323608 255134 323928 255218
rect 323608 254898 323650 255134
rect 323886 254898 323928 255134
rect 323608 254866 323928 254898
rect 354328 255454 354648 255486
rect 354328 255218 354370 255454
rect 354606 255218 354648 255454
rect 354328 255134 354648 255218
rect 354328 254898 354370 255134
rect 354606 254898 354648 255134
rect 354328 254866 354648 254898
rect 385048 255454 385368 255486
rect 385048 255218 385090 255454
rect 385326 255218 385368 255454
rect 385048 255134 385368 255218
rect 385048 254898 385090 255134
rect 385326 254898 385368 255134
rect 385048 254866 385368 254898
rect 415768 255454 416088 255486
rect 415768 255218 415810 255454
rect 416046 255218 416088 255454
rect 415768 255134 416088 255218
rect 415768 254898 415810 255134
rect 416046 254898 416088 255134
rect 415768 254866 416088 254898
rect 423234 244894 423854 280338
rect 423234 244658 423266 244894
rect 423502 244658 423586 244894
rect 423822 244658 423854 244894
rect 423234 244574 423854 244658
rect 423234 244338 423266 244574
rect 423502 244338 423586 244574
rect 423822 244338 423854 244574
rect 185368 237454 185688 237486
rect 185368 237218 185410 237454
rect 185646 237218 185688 237454
rect 185368 237134 185688 237218
rect 185368 236898 185410 237134
rect 185646 236898 185688 237134
rect 185368 236866 185688 236898
rect 216088 237454 216408 237486
rect 216088 237218 216130 237454
rect 216366 237218 216408 237454
rect 216088 237134 216408 237218
rect 216088 236898 216130 237134
rect 216366 236898 216408 237134
rect 216088 236866 216408 236898
rect 246808 237454 247128 237486
rect 246808 237218 246850 237454
rect 247086 237218 247128 237454
rect 246808 237134 247128 237218
rect 246808 236898 246850 237134
rect 247086 236898 247128 237134
rect 246808 236866 247128 236898
rect 277528 237454 277848 237486
rect 277528 237218 277570 237454
rect 277806 237218 277848 237454
rect 277528 237134 277848 237218
rect 277528 236898 277570 237134
rect 277806 236898 277848 237134
rect 277528 236866 277848 236898
rect 308248 237454 308568 237486
rect 308248 237218 308290 237454
rect 308526 237218 308568 237454
rect 308248 237134 308568 237218
rect 308248 236898 308290 237134
rect 308526 236898 308568 237134
rect 308248 236866 308568 236898
rect 338968 237454 339288 237486
rect 338968 237218 339010 237454
rect 339246 237218 339288 237454
rect 338968 237134 339288 237218
rect 338968 236898 339010 237134
rect 339246 236898 339288 237134
rect 338968 236866 339288 236898
rect 369688 237454 370008 237486
rect 369688 237218 369730 237454
rect 369966 237218 370008 237454
rect 369688 237134 370008 237218
rect 369688 236898 369730 237134
rect 369966 236898 370008 237134
rect 369688 236866 370008 236898
rect 400408 237454 400728 237486
rect 400408 237218 400450 237454
rect 400686 237218 400728 237454
rect 400408 237134 400728 237218
rect 400408 236898 400450 237134
rect 400686 236898 400728 237134
rect 400408 236866 400728 236898
rect 156954 230378 156986 230614
rect 157222 230378 157306 230614
rect 157542 230378 157574 230614
rect 156954 230294 157574 230378
rect 156954 230058 156986 230294
rect 157222 230058 157306 230294
rect 157542 230058 157574 230294
rect 156954 194614 157574 230058
rect 170008 219454 170328 219486
rect 170008 219218 170050 219454
rect 170286 219218 170328 219454
rect 170008 219134 170328 219218
rect 170008 218898 170050 219134
rect 170286 218898 170328 219134
rect 170008 218866 170328 218898
rect 200728 219454 201048 219486
rect 200728 219218 200770 219454
rect 201006 219218 201048 219454
rect 200728 219134 201048 219218
rect 200728 218898 200770 219134
rect 201006 218898 201048 219134
rect 200728 218866 201048 218898
rect 231448 219454 231768 219486
rect 231448 219218 231490 219454
rect 231726 219218 231768 219454
rect 231448 219134 231768 219218
rect 231448 218898 231490 219134
rect 231726 218898 231768 219134
rect 231448 218866 231768 218898
rect 262168 219454 262488 219486
rect 262168 219218 262210 219454
rect 262446 219218 262488 219454
rect 262168 219134 262488 219218
rect 262168 218898 262210 219134
rect 262446 218898 262488 219134
rect 262168 218866 262488 218898
rect 292888 219454 293208 219486
rect 292888 219218 292930 219454
rect 293166 219218 293208 219454
rect 292888 219134 293208 219218
rect 292888 218898 292930 219134
rect 293166 218898 293208 219134
rect 292888 218866 293208 218898
rect 323608 219454 323928 219486
rect 323608 219218 323650 219454
rect 323886 219218 323928 219454
rect 323608 219134 323928 219218
rect 323608 218898 323650 219134
rect 323886 218898 323928 219134
rect 323608 218866 323928 218898
rect 354328 219454 354648 219486
rect 354328 219218 354370 219454
rect 354606 219218 354648 219454
rect 354328 219134 354648 219218
rect 354328 218898 354370 219134
rect 354606 218898 354648 219134
rect 354328 218866 354648 218898
rect 385048 219454 385368 219486
rect 385048 219218 385090 219454
rect 385326 219218 385368 219454
rect 385048 219134 385368 219218
rect 385048 218898 385090 219134
rect 385326 218898 385368 219134
rect 385048 218866 385368 218898
rect 415768 219454 416088 219486
rect 415768 219218 415810 219454
rect 416046 219218 416088 219454
rect 415768 219134 416088 219218
rect 415768 218898 415810 219134
rect 416046 218898 416088 219134
rect 415768 218866 416088 218898
rect 423234 208894 423854 244338
rect 423234 208658 423266 208894
rect 423502 208658 423586 208894
rect 423822 208658 423854 208894
rect 423234 208574 423854 208658
rect 423234 208338 423266 208574
rect 423502 208338 423586 208574
rect 423822 208338 423854 208574
rect 156954 194378 156986 194614
rect 157222 194378 157306 194614
rect 157542 194378 157574 194614
rect 156954 194294 157574 194378
rect 156954 194058 156986 194294
rect 157222 194058 157306 194294
rect 157542 194058 157574 194294
rect 156954 158614 157574 194058
rect 156954 158378 156986 158614
rect 157222 158378 157306 158614
rect 157542 158378 157574 158614
rect 156954 158294 157574 158378
rect 156954 158058 156986 158294
rect 157222 158058 157306 158294
rect 157542 158058 157574 158294
rect 156954 122614 157574 158058
rect 156954 122378 156986 122614
rect 157222 122378 157306 122614
rect 157542 122378 157574 122614
rect 156954 122294 157574 122378
rect 156954 122058 156986 122294
rect 157222 122058 157306 122294
rect 157542 122058 157574 122294
rect 156954 86614 157574 122058
rect 156954 86378 156986 86614
rect 157222 86378 157306 86614
rect 157542 86378 157574 86614
rect 156954 86294 157574 86378
rect 156954 86058 156986 86294
rect 157222 86058 157306 86294
rect 157542 86058 157574 86294
rect 156954 50614 157574 86058
rect 156954 50378 156986 50614
rect 157222 50378 157306 50614
rect 157542 50378 157574 50614
rect 156954 50294 157574 50378
rect 156954 50058 156986 50294
rect 157222 50058 157306 50294
rect 157542 50058 157574 50294
rect 156954 14614 157574 50058
rect 156954 14378 156986 14614
rect 157222 14378 157306 14614
rect 157542 14378 157574 14614
rect 156954 14294 157574 14378
rect 156954 14058 156986 14294
rect 157222 14058 157306 14294
rect 157542 14058 157574 14294
rect 138954 -7302 138986 -7066
rect 139222 -7302 139306 -7066
rect 139542 -7302 139574 -7066
rect 138954 -7386 139574 -7302
rect 138954 -7622 138986 -7386
rect 139222 -7622 139306 -7386
rect 139542 -7622 139574 -7386
rect 138954 -7654 139574 -7622
rect 156954 -6106 157574 14058
rect 163794 165454 164414 198800
rect 163794 165218 163826 165454
rect 164062 165218 164146 165454
rect 164382 165218 164414 165454
rect 163794 165134 164414 165218
rect 163794 164898 163826 165134
rect 164062 164898 164146 165134
rect 164382 164898 164414 165134
rect 163794 129454 164414 164898
rect 163794 129218 163826 129454
rect 164062 129218 164146 129454
rect 164382 129218 164414 129454
rect 163794 129134 164414 129218
rect 163794 128898 163826 129134
rect 164062 128898 164146 129134
rect 164382 128898 164414 129134
rect 163794 93454 164414 128898
rect 163794 93218 163826 93454
rect 164062 93218 164146 93454
rect 164382 93218 164414 93454
rect 163794 93134 164414 93218
rect 163794 92898 163826 93134
rect 164062 92898 164146 93134
rect 164382 92898 164414 93134
rect 163794 57454 164414 92898
rect 163794 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 164414 57454
rect 163794 57134 164414 57218
rect 163794 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 164414 57134
rect 163794 21454 164414 56898
rect 163794 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 164414 21454
rect 163794 21134 164414 21218
rect 163794 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 164414 21134
rect 163794 -1306 164414 20898
rect 163794 -1542 163826 -1306
rect 164062 -1542 164146 -1306
rect 164382 -1542 164414 -1306
rect 163794 -1626 164414 -1542
rect 163794 -1862 163826 -1626
rect 164062 -1862 164146 -1626
rect 164382 -1862 164414 -1626
rect 163794 -1894 164414 -1862
rect 167514 169174 168134 198800
rect 167514 168938 167546 169174
rect 167782 168938 167866 169174
rect 168102 168938 168134 169174
rect 167514 168854 168134 168938
rect 167514 168618 167546 168854
rect 167782 168618 167866 168854
rect 168102 168618 168134 168854
rect 167514 133174 168134 168618
rect 167514 132938 167546 133174
rect 167782 132938 167866 133174
rect 168102 132938 168134 133174
rect 167514 132854 168134 132938
rect 167514 132618 167546 132854
rect 167782 132618 167866 132854
rect 168102 132618 168134 132854
rect 167514 97174 168134 132618
rect 167514 96938 167546 97174
rect 167782 96938 167866 97174
rect 168102 96938 168134 97174
rect 167514 96854 168134 96938
rect 167514 96618 167546 96854
rect 167782 96618 167866 96854
rect 168102 96618 168134 96854
rect 167514 61174 168134 96618
rect 167514 60938 167546 61174
rect 167782 60938 167866 61174
rect 168102 60938 168134 61174
rect 167514 60854 168134 60938
rect 167514 60618 167546 60854
rect 167782 60618 167866 60854
rect 168102 60618 168134 60854
rect 167514 25174 168134 60618
rect 167514 24938 167546 25174
rect 167782 24938 167866 25174
rect 168102 24938 168134 25174
rect 167514 24854 168134 24938
rect 167514 24618 167546 24854
rect 167782 24618 167866 24854
rect 168102 24618 168134 24854
rect 167514 -3226 168134 24618
rect 167514 -3462 167546 -3226
rect 167782 -3462 167866 -3226
rect 168102 -3462 168134 -3226
rect 167514 -3546 168134 -3462
rect 167514 -3782 167546 -3546
rect 167782 -3782 167866 -3546
rect 168102 -3782 168134 -3546
rect 167514 -3814 168134 -3782
rect 171234 172894 171854 198800
rect 171234 172658 171266 172894
rect 171502 172658 171586 172894
rect 171822 172658 171854 172894
rect 171234 172574 171854 172658
rect 171234 172338 171266 172574
rect 171502 172338 171586 172574
rect 171822 172338 171854 172574
rect 171234 136894 171854 172338
rect 171234 136658 171266 136894
rect 171502 136658 171586 136894
rect 171822 136658 171854 136894
rect 171234 136574 171854 136658
rect 171234 136338 171266 136574
rect 171502 136338 171586 136574
rect 171822 136338 171854 136574
rect 171234 100894 171854 136338
rect 171234 100658 171266 100894
rect 171502 100658 171586 100894
rect 171822 100658 171854 100894
rect 171234 100574 171854 100658
rect 171234 100338 171266 100574
rect 171502 100338 171586 100574
rect 171822 100338 171854 100574
rect 171234 64894 171854 100338
rect 171234 64658 171266 64894
rect 171502 64658 171586 64894
rect 171822 64658 171854 64894
rect 171234 64574 171854 64658
rect 171234 64338 171266 64574
rect 171502 64338 171586 64574
rect 171822 64338 171854 64574
rect 171234 28894 171854 64338
rect 171234 28658 171266 28894
rect 171502 28658 171586 28894
rect 171822 28658 171854 28894
rect 171234 28574 171854 28658
rect 171234 28338 171266 28574
rect 171502 28338 171586 28574
rect 171822 28338 171854 28574
rect 171234 -5146 171854 28338
rect 171234 -5382 171266 -5146
rect 171502 -5382 171586 -5146
rect 171822 -5382 171854 -5146
rect 171234 -5466 171854 -5382
rect 171234 -5702 171266 -5466
rect 171502 -5702 171586 -5466
rect 171822 -5702 171854 -5466
rect 171234 -5734 171854 -5702
rect 174954 176614 175574 198800
rect 174954 176378 174986 176614
rect 175222 176378 175306 176614
rect 175542 176378 175574 176614
rect 174954 176294 175574 176378
rect 174954 176058 174986 176294
rect 175222 176058 175306 176294
rect 175542 176058 175574 176294
rect 174954 140614 175574 176058
rect 174954 140378 174986 140614
rect 175222 140378 175306 140614
rect 175542 140378 175574 140614
rect 174954 140294 175574 140378
rect 174954 140058 174986 140294
rect 175222 140058 175306 140294
rect 175542 140058 175574 140294
rect 174954 104614 175574 140058
rect 174954 104378 174986 104614
rect 175222 104378 175306 104614
rect 175542 104378 175574 104614
rect 174954 104294 175574 104378
rect 174954 104058 174986 104294
rect 175222 104058 175306 104294
rect 175542 104058 175574 104294
rect 174954 68614 175574 104058
rect 174954 68378 174986 68614
rect 175222 68378 175306 68614
rect 175542 68378 175574 68614
rect 174954 68294 175574 68378
rect 174954 68058 174986 68294
rect 175222 68058 175306 68294
rect 175542 68058 175574 68294
rect 174954 32614 175574 68058
rect 174954 32378 174986 32614
rect 175222 32378 175306 32614
rect 175542 32378 175574 32614
rect 174954 32294 175574 32378
rect 174954 32058 174986 32294
rect 175222 32058 175306 32294
rect 175542 32058 175574 32294
rect 156954 -6342 156986 -6106
rect 157222 -6342 157306 -6106
rect 157542 -6342 157574 -6106
rect 156954 -6426 157574 -6342
rect 156954 -6662 156986 -6426
rect 157222 -6662 157306 -6426
rect 157542 -6662 157574 -6426
rect 156954 -7654 157574 -6662
rect 174954 -7066 175574 32058
rect 181794 183454 182414 198800
rect 181794 183218 181826 183454
rect 182062 183218 182146 183454
rect 182382 183218 182414 183454
rect 181794 183134 182414 183218
rect 181794 182898 181826 183134
rect 182062 182898 182146 183134
rect 182382 182898 182414 183134
rect 181794 147454 182414 182898
rect 181794 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 182414 147454
rect 181794 147134 182414 147218
rect 181794 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 182414 147134
rect 181794 111454 182414 146898
rect 181794 111218 181826 111454
rect 182062 111218 182146 111454
rect 182382 111218 182414 111454
rect 181794 111134 182414 111218
rect 181794 110898 181826 111134
rect 182062 110898 182146 111134
rect 182382 110898 182414 111134
rect 181794 75454 182414 110898
rect 181794 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 182414 75454
rect 181794 75134 182414 75218
rect 181794 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 182414 75134
rect 181794 39454 182414 74898
rect 181794 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 182414 39454
rect 181794 39134 182414 39218
rect 181794 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 182414 39134
rect 181794 3454 182414 38898
rect 181794 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 182414 3454
rect 181794 3134 182414 3218
rect 181794 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 182414 3134
rect 181794 -346 182414 2898
rect 181794 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 182414 -346
rect 181794 -666 182414 -582
rect 181794 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 182414 -666
rect 181794 -1894 182414 -902
rect 185514 187174 186134 198800
rect 185514 186938 185546 187174
rect 185782 186938 185866 187174
rect 186102 186938 186134 187174
rect 185514 186854 186134 186938
rect 185514 186618 185546 186854
rect 185782 186618 185866 186854
rect 186102 186618 186134 186854
rect 185514 151174 186134 186618
rect 185514 150938 185546 151174
rect 185782 150938 185866 151174
rect 186102 150938 186134 151174
rect 185514 150854 186134 150938
rect 185514 150618 185546 150854
rect 185782 150618 185866 150854
rect 186102 150618 186134 150854
rect 185514 115174 186134 150618
rect 185514 114938 185546 115174
rect 185782 114938 185866 115174
rect 186102 114938 186134 115174
rect 185514 114854 186134 114938
rect 185514 114618 185546 114854
rect 185782 114618 185866 114854
rect 186102 114618 186134 114854
rect 185514 79174 186134 114618
rect 185514 78938 185546 79174
rect 185782 78938 185866 79174
rect 186102 78938 186134 79174
rect 185514 78854 186134 78938
rect 185514 78618 185546 78854
rect 185782 78618 185866 78854
rect 186102 78618 186134 78854
rect 185514 43174 186134 78618
rect 185514 42938 185546 43174
rect 185782 42938 185866 43174
rect 186102 42938 186134 43174
rect 185514 42854 186134 42938
rect 185514 42618 185546 42854
rect 185782 42618 185866 42854
rect 186102 42618 186134 42854
rect 185514 7174 186134 42618
rect 185514 6938 185546 7174
rect 185782 6938 185866 7174
rect 186102 6938 186134 7174
rect 185514 6854 186134 6938
rect 185514 6618 185546 6854
rect 185782 6618 185866 6854
rect 186102 6618 186134 6854
rect 185514 -2266 186134 6618
rect 185514 -2502 185546 -2266
rect 185782 -2502 185866 -2266
rect 186102 -2502 186134 -2266
rect 185514 -2586 186134 -2502
rect 185514 -2822 185546 -2586
rect 185782 -2822 185866 -2586
rect 186102 -2822 186134 -2586
rect 185514 -3814 186134 -2822
rect 189234 190894 189854 198800
rect 189234 190658 189266 190894
rect 189502 190658 189586 190894
rect 189822 190658 189854 190894
rect 189234 190574 189854 190658
rect 189234 190338 189266 190574
rect 189502 190338 189586 190574
rect 189822 190338 189854 190574
rect 189234 154894 189854 190338
rect 189234 154658 189266 154894
rect 189502 154658 189586 154894
rect 189822 154658 189854 154894
rect 189234 154574 189854 154658
rect 189234 154338 189266 154574
rect 189502 154338 189586 154574
rect 189822 154338 189854 154574
rect 189234 118894 189854 154338
rect 189234 118658 189266 118894
rect 189502 118658 189586 118894
rect 189822 118658 189854 118894
rect 189234 118574 189854 118658
rect 189234 118338 189266 118574
rect 189502 118338 189586 118574
rect 189822 118338 189854 118574
rect 189234 82894 189854 118338
rect 189234 82658 189266 82894
rect 189502 82658 189586 82894
rect 189822 82658 189854 82894
rect 189234 82574 189854 82658
rect 189234 82338 189266 82574
rect 189502 82338 189586 82574
rect 189822 82338 189854 82574
rect 189234 46894 189854 82338
rect 189234 46658 189266 46894
rect 189502 46658 189586 46894
rect 189822 46658 189854 46894
rect 189234 46574 189854 46658
rect 189234 46338 189266 46574
rect 189502 46338 189586 46574
rect 189822 46338 189854 46574
rect 189234 10894 189854 46338
rect 189234 10658 189266 10894
rect 189502 10658 189586 10894
rect 189822 10658 189854 10894
rect 189234 10574 189854 10658
rect 189234 10338 189266 10574
rect 189502 10338 189586 10574
rect 189822 10338 189854 10574
rect 189234 -4186 189854 10338
rect 189234 -4422 189266 -4186
rect 189502 -4422 189586 -4186
rect 189822 -4422 189854 -4186
rect 189234 -4506 189854 -4422
rect 189234 -4742 189266 -4506
rect 189502 -4742 189586 -4506
rect 189822 -4742 189854 -4506
rect 189234 -5734 189854 -4742
rect 192954 194614 193574 198800
rect 192954 194378 192986 194614
rect 193222 194378 193306 194614
rect 193542 194378 193574 194614
rect 192954 194294 193574 194378
rect 192954 194058 192986 194294
rect 193222 194058 193306 194294
rect 193542 194058 193574 194294
rect 192954 158614 193574 194058
rect 192954 158378 192986 158614
rect 193222 158378 193306 158614
rect 193542 158378 193574 158614
rect 192954 158294 193574 158378
rect 192954 158058 192986 158294
rect 193222 158058 193306 158294
rect 193542 158058 193574 158294
rect 192954 122614 193574 158058
rect 192954 122378 192986 122614
rect 193222 122378 193306 122614
rect 193542 122378 193574 122614
rect 192954 122294 193574 122378
rect 192954 122058 192986 122294
rect 193222 122058 193306 122294
rect 193542 122058 193574 122294
rect 192954 86614 193574 122058
rect 192954 86378 192986 86614
rect 193222 86378 193306 86614
rect 193542 86378 193574 86614
rect 192954 86294 193574 86378
rect 192954 86058 192986 86294
rect 193222 86058 193306 86294
rect 193542 86058 193574 86294
rect 192954 50614 193574 86058
rect 192954 50378 192986 50614
rect 193222 50378 193306 50614
rect 193542 50378 193574 50614
rect 192954 50294 193574 50378
rect 192954 50058 192986 50294
rect 193222 50058 193306 50294
rect 193542 50058 193574 50294
rect 192954 14614 193574 50058
rect 192954 14378 192986 14614
rect 193222 14378 193306 14614
rect 193542 14378 193574 14614
rect 192954 14294 193574 14378
rect 192954 14058 192986 14294
rect 193222 14058 193306 14294
rect 193542 14058 193574 14294
rect 174954 -7302 174986 -7066
rect 175222 -7302 175306 -7066
rect 175542 -7302 175574 -7066
rect 174954 -7386 175574 -7302
rect 174954 -7622 174986 -7386
rect 175222 -7622 175306 -7386
rect 175542 -7622 175574 -7386
rect 174954 -7654 175574 -7622
rect 192954 -6106 193574 14058
rect 199794 165454 200414 198800
rect 199794 165218 199826 165454
rect 200062 165218 200146 165454
rect 200382 165218 200414 165454
rect 199794 165134 200414 165218
rect 199794 164898 199826 165134
rect 200062 164898 200146 165134
rect 200382 164898 200414 165134
rect 199794 129454 200414 164898
rect 199794 129218 199826 129454
rect 200062 129218 200146 129454
rect 200382 129218 200414 129454
rect 199794 129134 200414 129218
rect 199794 128898 199826 129134
rect 200062 128898 200146 129134
rect 200382 128898 200414 129134
rect 199794 93454 200414 128898
rect 199794 93218 199826 93454
rect 200062 93218 200146 93454
rect 200382 93218 200414 93454
rect 199794 93134 200414 93218
rect 199794 92898 199826 93134
rect 200062 92898 200146 93134
rect 200382 92898 200414 93134
rect 199794 57454 200414 92898
rect 199794 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 200414 57454
rect 199794 57134 200414 57218
rect 199794 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 200414 57134
rect 199794 21454 200414 56898
rect 199794 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 200414 21454
rect 199794 21134 200414 21218
rect 199794 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 200414 21134
rect 199794 -1306 200414 20898
rect 199794 -1542 199826 -1306
rect 200062 -1542 200146 -1306
rect 200382 -1542 200414 -1306
rect 199794 -1626 200414 -1542
rect 199794 -1862 199826 -1626
rect 200062 -1862 200146 -1626
rect 200382 -1862 200414 -1626
rect 199794 -1894 200414 -1862
rect 203514 169174 204134 198800
rect 203514 168938 203546 169174
rect 203782 168938 203866 169174
rect 204102 168938 204134 169174
rect 203514 168854 204134 168938
rect 203514 168618 203546 168854
rect 203782 168618 203866 168854
rect 204102 168618 204134 168854
rect 203514 133174 204134 168618
rect 203514 132938 203546 133174
rect 203782 132938 203866 133174
rect 204102 132938 204134 133174
rect 203514 132854 204134 132938
rect 203514 132618 203546 132854
rect 203782 132618 203866 132854
rect 204102 132618 204134 132854
rect 203514 97174 204134 132618
rect 203514 96938 203546 97174
rect 203782 96938 203866 97174
rect 204102 96938 204134 97174
rect 203514 96854 204134 96938
rect 203514 96618 203546 96854
rect 203782 96618 203866 96854
rect 204102 96618 204134 96854
rect 203514 61174 204134 96618
rect 203514 60938 203546 61174
rect 203782 60938 203866 61174
rect 204102 60938 204134 61174
rect 203514 60854 204134 60938
rect 203514 60618 203546 60854
rect 203782 60618 203866 60854
rect 204102 60618 204134 60854
rect 203514 25174 204134 60618
rect 203514 24938 203546 25174
rect 203782 24938 203866 25174
rect 204102 24938 204134 25174
rect 203514 24854 204134 24938
rect 203514 24618 203546 24854
rect 203782 24618 203866 24854
rect 204102 24618 204134 24854
rect 203514 -3226 204134 24618
rect 203514 -3462 203546 -3226
rect 203782 -3462 203866 -3226
rect 204102 -3462 204134 -3226
rect 203514 -3546 204134 -3462
rect 203514 -3782 203546 -3546
rect 203782 -3782 203866 -3546
rect 204102 -3782 204134 -3546
rect 203514 -3814 204134 -3782
rect 207234 172894 207854 198800
rect 207234 172658 207266 172894
rect 207502 172658 207586 172894
rect 207822 172658 207854 172894
rect 207234 172574 207854 172658
rect 207234 172338 207266 172574
rect 207502 172338 207586 172574
rect 207822 172338 207854 172574
rect 207234 136894 207854 172338
rect 207234 136658 207266 136894
rect 207502 136658 207586 136894
rect 207822 136658 207854 136894
rect 207234 136574 207854 136658
rect 207234 136338 207266 136574
rect 207502 136338 207586 136574
rect 207822 136338 207854 136574
rect 207234 100894 207854 136338
rect 207234 100658 207266 100894
rect 207502 100658 207586 100894
rect 207822 100658 207854 100894
rect 207234 100574 207854 100658
rect 207234 100338 207266 100574
rect 207502 100338 207586 100574
rect 207822 100338 207854 100574
rect 207234 64894 207854 100338
rect 207234 64658 207266 64894
rect 207502 64658 207586 64894
rect 207822 64658 207854 64894
rect 207234 64574 207854 64658
rect 207234 64338 207266 64574
rect 207502 64338 207586 64574
rect 207822 64338 207854 64574
rect 207234 28894 207854 64338
rect 207234 28658 207266 28894
rect 207502 28658 207586 28894
rect 207822 28658 207854 28894
rect 207234 28574 207854 28658
rect 207234 28338 207266 28574
rect 207502 28338 207586 28574
rect 207822 28338 207854 28574
rect 207234 -5146 207854 28338
rect 207234 -5382 207266 -5146
rect 207502 -5382 207586 -5146
rect 207822 -5382 207854 -5146
rect 207234 -5466 207854 -5382
rect 207234 -5702 207266 -5466
rect 207502 -5702 207586 -5466
rect 207822 -5702 207854 -5466
rect 207234 -5734 207854 -5702
rect 210954 176614 211574 198800
rect 210954 176378 210986 176614
rect 211222 176378 211306 176614
rect 211542 176378 211574 176614
rect 210954 176294 211574 176378
rect 210954 176058 210986 176294
rect 211222 176058 211306 176294
rect 211542 176058 211574 176294
rect 210954 140614 211574 176058
rect 210954 140378 210986 140614
rect 211222 140378 211306 140614
rect 211542 140378 211574 140614
rect 210954 140294 211574 140378
rect 210954 140058 210986 140294
rect 211222 140058 211306 140294
rect 211542 140058 211574 140294
rect 210954 104614 211574 140058
rect 210954 104378 210986 104614
rect 211222 104378 211306 104614
rect 211542 104378 211574 104614
rect 210954 104294 211574 104378
rect 210954 104058 210986 104294
rect 211222 104058 211306 104294
rect 211542 104058 211574 104294
rect 210954 68614 211574 104058
rect 210954 68378 210986 68614
rect 211222 68378 211306 68614
rect 211542 68378 211574 68614
rect 210954 68294 211574 68378
rect 210954 68058 210986 68294
rect 211222 68058 211306 68294
rect 211542 68058 211574 68294
rect 210954 32614 211574 68058
rect 210954 32378 210986 32614
rect 211222 32378 211306 32614
rect 211542 32378 211574 32614
rect 210954 32294 211574 32378
rect 210954 32058 210986 32294
rect 211222 32058 211306 32294
rect 211542 32058 211574 32294
rect 192954 -6342 192986 -6106
rect 193222 -6342 193306 -6106
rect 193542 -6342 193574 -6106
rect 192954 -6426 193574 -6342
rect 192954 -6662 192986 -6426
rect 193222 -6662 193306 -6426
rect 193542 -6662 193574 -6426
rect 192954 -7654 193574 -6662
rect 210954 -7066 211574 32058
rect 217794 183454 218414 198800
rect 217794 183218 217826 183454
rect 218062 183218 218146 183454
rect 218382 183218 218414 183454
rect 217794 183134 218414 183218
rect 217794 182898 217826 183134
rect 218062 182898 218146 183134
rect 218382 182898 218414 183134
rect 217794 147454 218414 182898
rect 217794 147218 217826 147454
rect 218062 147218 218146 147454
rect 218382 147218 218414 147454
rect 217794 147134 218414 147218
rect 217794 146898 217826 147134
rect 218062 146898 218146 147134
rect 218382 146898 218414 147134
rect 217794 111454 218414 146898
rect 217794 111218 217826 111454
rect 218062 111218 218146 111454
rect 218382 111218 218414 111454
rect 217794 111134 218414 111218
rect 217794 110898 217826 111134
rect 218062 110898 218146 111134
rect 218382 110898 218414 111134
rect 217794 75454 218414 110898
rect 217794 75218 217826 75454
rect 218062 75218 218146 75454
rect 218382 75218 218414 75454
rect 217794 75134 218414 75218
rect 217794 74898 217826 75134
rect 218062 74898 218146 75134
rect 218382 74898 218414 75134
rect 217794 39454 218414 74898
rect 217794 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 218414 39454
rect 217794 39134 218414 39218
rect 217794 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 218414 39134
rect 217794 3454 218414 38898
rect 217794 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 218414 3454
rect 217794 3134 218414 3218
rect 217794 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 218414 3134
rect 217794 -346 218414 2898
rect 217794 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 218414 -346
rect 217794 -666 218414 -582
rect 217794 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 218414 -666
rect 217794 -1894 218414 -902
rect 221514 187174 222134 198800
rect 221514 186938 221546 187174
rect 221782 186938 221866 187174
rect 222102 186938 222134 187174
rect 221514 186854 222134 186938
rect 221514 186618 221546 186854
rect 221782 186618 221866 186854
rect 222102 186618 222134 186854
rect 221514 151174 222134 186618
rect 221514 150938 221546 151174
rect 221782 150938 221866 151174
rect 222102 150938 222134 151174
rect 221514 150854 222134 150938
rect 221514 150618 221546 150854
rect 221782 150618 221866 150854
rect 222102 150618 222134 150854
rect 221514 115174 222134 150618
rect 221514 114938 221546 115174
rect 221782 114938 221866 115174
rect 222102 114938 222134 115174
rect 221514 114854 222134 114938
rect 221514 114618 221546 114854
rect 221782 114618 221866 114854
rect 222102 114618 222134 114854
rect 221514 79174 222134 114618
rect 221514 78938 221546 79174
rect 221782 78938 221866 79174
rect 222102 78938 222134 79174
rect 221514 78854 222134 78938
rect 221514 78618 221546 78854
rect 221782 78618 221866 78854
rect 222102 78618 222134 78854
rect 221514 43174 222134 78618
rect 221514 42938 221546 43174
rect 221782 42938 221866 43174
rect 222102 42938 222134 43174
rect 221514 42854 222134 42938
rect 221514 42618 221546 42854
rect 221782 42618 221866 42854
rect 222102 42618 222134 42854
rect 221514 7174 222134 42618
rect 221514 6938 221546 7174
rect 221782 6938 221866 7174
rect 222102 6938 222134 7174
rect 221514 6854 222134 6938
rect 221514 6618 221546 6854
rect 221782 6618 221866 6854
rect 222102 6618 222134 6854
rect 221514 -2266 222134 6618
rect 221514 -2502 221546 -2266
rect 221782 -2502 221866 -2266
rect 222102 -2502 222134 -2266
rect 221514 -2586 222134 -2502
rect 221514 -2822 221546 -2586
rect 221782 -2822 221866 -2586
rect 222102 -2822 222134 -2586
rect 221514 -3814 222134 -2822
rect 225234 190894 225854 198800
rect 225234 190658 225266 190894
rect 225502 190658 225586 190894
rect 225822 190658 225854 190894
rect 225234 190574 225854 190658
rect 225234 190338 225266 190574
rect 225502 190338 225586 190574
rect 225822 190338 225854 190574
rect 225234 154894 225854 190338
rect 225234 154658 225266 154894
rect 225502 154658 225586 154894
rect 225822 154658 225854 154894
rect 225234 154574 225854 154658
rect 225234 154338 225266 154574
rect 225502 154338 225586 154574
rect 225822 154338 225854 154574
rect 225234 118894 225854 154338
rect 225234 118658 225266 118894
rect 225502 118658 225586 118894
rect 225822 118658 225854 118894
rect 225234 118574 225854 118658
rect 225234 118338 225266 118574
rect 225502 118338 225586 118574
rect 225822 118338 225854 118574
rect 225234 82894 225854 118338
rect 225234 82658 225266 82894
rect 225502 82658 225586 82894
rect 225822 82658 225854 82894
rect 225234 82574 225854 82658
rect 225234 82338 225266 82574
rect 225502 82338 225586 82574
rect 225822 82338 225854 82574
rect 225234 46894 225854 82338
rect 225234 46658 225266 46894
rect 225502 46658 225586 46894
rect 225822 46658 225854 46894
rect 225234 46574 225854 46658
rect 225234 46338 225266 46574
rect 225502 46338 225586 46574
rect 225822 46338 225854 46574
rect 225234 10894 225854 46338
rect 225234 10658 225266 10894
rect 225502 10658 225586 10894
rect 225822 10658 225854 10894
rect 225234 10574 225854 10658
rect 225234 10338 225266 10574
rect 225502 10338 225586 10574
rect 225822 10338 225854 10574
rect 225234 -4186 225854 10338
rect 225234 -4422 225266 -4186
rect 225502 -4422 225586 -4186
rect 225822 -4422 225854 -4186
rect 225234 -4506 225854 -4422
rect 225234 -4742 225266 -4506
rect 225502 -4742 225586 -4506
rect 225822 -4742 225854 -4506
rect 225234 -5734 225854 -4742
rect 228954 194614 229574 198800
rect 228954 194378 228986 194614
rect 229222 194378 229306 194614
rect 229542 194378 229574 194614
rect 228954 194294 229574 194378
rect 228954 194058 228986 194294
rect 229222 194058 229306 194294
rect 229542 194058 229574 194294
rect 228954 158614 229574 194058
rect 228954 158378 228986 158614
rect 229222 158378 229306 158614
rect 229542 158378 229574 158614
rect 228954 158294 229574 158378
rect 228954 158058 228986 158294
rect 229222 158058 229306 158294
rect 229542 158058 229574 158294
rect 228954 122614 229574 158058
rect 228954 122378 228986 122614
rect 229222 122378 229306 122614
rect 229542 122378 229574 122614
rect 228954 122294 229574 122378
rect 228954 122058 228986 122294
rect 229222 122058 229306 122294
rect 229542 122058 229574 122294
rect 228954 86614 229574 122058
rect 228954 86378 228986 86614
rect 229222 86378 229306 86614
rect 229542 86378 229574 86614
rect 228954 86294 229574 86378
rect 228954 86058 228986 86294
rect 229222 86058 229306 86294
rect 229542 86058 229574 86294
rect 228954 50614 229574 86058
rect 228954 50378 228986 50614
rect 229222 50378 229306 50614
rect 229542 50378 229574 50614
rect 228954 50294 229574 50378
rect 228954 50058 228986 50294
rect 229222 50058 229306 50294
rect 229542 50058 229574 50294
rect 228954 14614 229574 50058
rect 228954 14378 228986 14614
rect 229222 14378 229306 14614
rect 229542 14378 229574 14614
rect 228954 14294 229574 14378
rect 228954 14058 228986 14294
rect 229222 14058 229306 14294
rect 229542 14058 229574 14294
rect 210954 -7302 210986 -7066
rect 211222 -7302 211306 -7066
rect 211542 -7302 211574 -7066
rect 210954 -7386 211574 -7302
rect 210954 -7622 210986 -7386
rect 211222 -7622 211306 -7386
rect 211542 -7622 211574 -7386
rect 210954 -7654 211574 -7622
rect 228954 -6106 229574 14058
rect 235794 165454 236414 198800
rect 235794 165218 235826 165454
rect 236062 165218 236146 165454
rect 236382 165218 236414 165454
rect 235794 165134 236414 165218
rect 235794 164898 235826 165134
rect 236062 164898 236146 165134
rect 236382 164898 236414 165134
rect 235794 129454 236414 164898
rect 235794 129218 235826 129454
rect 236062 129218 236146 129454
rect 236382 129218 236414 129454
rect 235794 129134 236414 129218
rect 235794 128898 235826 129134
rect 236062 128898 236146 129134
rect 236382 128898 236414 129134
rect 235794 93454 236414 128898
rect 235794 93218 235826 93454
rect 236062 93218 236146 93454
rect 236382 93218 236414 93454
rect 235794 93134 236414 93218
rect 235794 92898 235826 93134
rect 236062 92898 236146 93134
rect 236382 92898 236414 93134
rect 235794 57454 236414 92898
rect 235794 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 236414 57454
rect 235794 57134 236414 57218
rect 235794 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 236414 57134
rect 235794 21454 236414 56898
rect 235794 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 236414 21454
rect 235794 21134 236414 21218
rect 235794 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 236414 21134
rect 235794 -1306 236414 20898
rect 235794 -1542 235826 -1306
rect 236062 -1542 236146 -1306
rect 236382 -1542 236414 -1306
rect 235794 -1626 236414 -1542
rect 235794 -1862 235826 -1626
rect 236062 -1862 236146 -1626
rect 236382 -1862 236414 -1626
rect 235794 -1894 236414 -1862
rect 239514 169174 240134 198800
rect 239514 168938 239546 169174
rect 239782 168938 239866 169174
rect 240102 168938 240134 169174
rect 239514 168854 240134 168938
rect 239514 168618 239546 168854
rect 239782 168618 239866 168854
rect 240102 168618 240134 168854
rect 239514 133174 240134 168618
rect 239514 132938 239546 133174
rect 239782 132938 239866 133174
rect 240102 132938 240134 133174
rect 239514 132854 240134 132938
rect 239514 132618 239546 132854
rect 239782 132618 239866 132854
rect 240102 132618 240134 132854
rect 239514 97174 240134 132618
rect 239514 96938 239546 97174
rect 239782 96938 239866 97174
rect 240102 96938 240134 97174
rect 239514 96854 240134 96938
rect 239514 96618 239546 96854
rect 239782 96618 239866 96854
rect 240102 96618 240134 96854
rect 239514 61174 240134 96618
rect 239514 60938 239546 61174
rect 239782 60938 239866 61174
rect 240102 60938 240134 61174
rect 239514 60854 240134 60938
rect 239514 60618 239546 60854
rect 239782 60618 239866 60854
rect 240102 60618 240134 60854
rect 239514 25174 240134 60618
rect 239514 24938 239546 25174
rect 239782 24938 239866 25174
rect 240102 24938 240134 25174
rect 239514 24854 240134 24938
rect 239514 24618 239546 24854
rect 239782 24618 239866 24854
rect 240102 24618 240134 24854
rect 239514 -3226 240134 24618
rect 239514 -3462 239546 -3226
rect 239782 -3462 239866 -3226
rect 240102 -3462 240134 -3226
rect 239514 -3546 240134 -3462
rect 239514 -3782 239546 -3546
rect 239782 -3782 239866 -3546
rect 240102 -3782 240134 -3546
rect 239514 -3814 240134 -3782
rect 243234 172894 243854 198800
rect 243234 172658 243266 172894
rect 243502 172658 243586 172894
rect 243822 172658 243854 172894
rect 243234 172574 243854 172658
rect 243234 172338 243266 172574
rect 243502 172338 243586 172574
rect 243822 172338 243854 172574
rect 243234 136894 243854 172338
rect 243234 136658 243266 136894
rect 243502 136658 243586 136894
rect 243822 136658 243854 136894
rect 243234 136574 243854 136658
rect 243234 136338 243266 136574
rect 243502 136338 243586 136574
rect 243822 136338 243854 136574
rect 243234 100894 243854 136338
rect 243234 100658 243266 100894
rect 243502 100658 243586 100894
rect 243822 100658 243854 100894
rect 243234 100574 243854 100658
rect 243234 100338 243266 100574
rect 243502 100338 243586 100574
rect 243822 100338 243854 100574
rect 243234 64894 243854 100338
rect 243234 64658 243266 64894
rect 243502 64658 243586 64894
rect 243822 64658 243854 64894
rect 243234 64574 243854 64658
rect 243234 64338 243266 64574
rect 243502 64338 243586 64574
rect 243822 64338 243854 64574
rect 243234 28894 243854 64338
rect 243234 28658 243266 28894
rect 243502 28658 243586 28894
rect 243822 28658 243854 28894
rect 243234 28574 243854 28658
rect 243234 28338 243266 28574
rect 243502 28338 243586 28574
rect 243822 28338 243854 28574
rect 243234 -5146 243854 28338
rect 243234 -5382 243266 -5146
rect 243502 -5382 243586 -5146
rect 243822 -5382 243854 -5146
rect 243234 -5466 243854 -5382
rect 243234 -5702 243266 -5466
rect 243502 -5702 243586 -5466
rect 243822 -5702 243854 -5466
rect 243234 -5734 243854 -5702
rect 246954 176614 247574 198800
rect 246954 176378 246986 176614
rect 247222 176378 247306 176614
rect 247542 176378 247574 176614
rect 246954 176294 247574 176378
rect 246954 176058 246986 176294
rect 247222 176058 247306 176294
rect 247542 176058 247574 176294
rect 246954 140614 247574 176058
rect 246954 140378 246986 140614
rect 247222 140378 247306 140614
rect 247542 140378 247574 140614
rect 246954 140294 247574 140378
rect 246954 140058 246986 140294
rect 247222 140058 247306 140294
rect 247542 140058 247574 140294
rect 246954 104614 247574 140058
rect 246954 104378 246986 104614
rect 247222 104378 247306 104614
rect 247542 104378 247574 104614
rect 246954 104294 247574 104378
rect 246954 104058 246986 104294
rect 247222 104058 247306 104294
rect 247542 104058 247574 104294
rect 246954 68614 247574 104058
rect 246954 68378 246986 68614
rect 247222 68378 247306 68614
rect 247542 68378 247574 68614
rect 246954 68294 247574 68378
rect 246954 68058 246986 68294
rect 247222 68058 247306 68294
rect 247542 68058 247574 68294
rect 246954 32614 247574 68058
rect 246954 32378 246986 32614
rect 247222 32378 247306 32614
rect 247542 32378 247574 32614
rect 246954 32294 247574 32378
rect 246954 32058 246986 32294
rect 247222 32058 247306 32294
rect 247542 32058 247574 32294
rect 228954 -6342 228986 -6106
rect 229222 -6342 229306 -6106
rect 229542 -6342 229574 -6106
rect 228954 -6426 229574 -6342
rect 228954 -6662 228986 -6426
rect 229222 -6662 229306 -6426
rect 229542 -6662 229574 -6426
rect 228954 -7654 229574 -6662
rect 246954 -7066 247574 32058
rect 253794 183454 254414 198800
rect 253794 183218 253826 183454
rect 254062 183218 254146 183454
rect 254382 183218 254414 183454
rect 253794 183134 254414 183218
rect 253794 182898 253826 183134
rect 254062 182898 254146 183134
rect 254382 182898 254414 183134
rect 253794 147454 254414 182898
rect 253794 147218 253826 147454
rect 254062 147218 254146 147454
rect 254382 147218 254414 147454
rect 253794 147134 254414 147218
rect 253794 146898 253826 147134
rect 254062 146898 254146 147134
rect 254382 146898 254414 147134
rect 253794 111454 254414 146898
rect 253794 111218 253826 111454
rect 254062 111218 254146 111454
rect 254382 111218 254414 111454
rect 253794 111134 254414 111218
rect 253794 110898 253826 111134
rect 254062 110898 254146 111134
rect 254382 110898 254414 111134
rect 253794 75454 254414 110898
rect 253794 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 254414 75454
rect 253794 75134 254414 75218
rect 253794 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 254414 75134
rect 253794 39454 254414 74898
rect 253794 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 254414 39454
rect 253794 39134 254414 39218
rect 253794 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 254414 39134
rect 253794 3454 254414 38898
rect 253794 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 254414 3454
rect 253794 3134 254414 3218
rect 253794 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 254414 3134
rect 253794 -346 254414 2898
rect 253794 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 254414 -346
rect 253794 -666 254414 -582
rect 253794 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 254414 -666
rect 253794 -1894 254414 -902
rect 257514 187174 258134 198800
rect 257514 186938 257546 187174
rect 257782 186938 257866 187174
rect 258102 186938 258134 187174
rect 257514 186854 258134 186938
rect 257514 186618 257546 186854
rect 257782 186618 257866 186854
rect 258102 186618 258134 186854
rect 257514 151174 258134 186618
rect 257514 150938 257546 151174
rect 257782 150938 257866 151174
rect 258102 150938 258134 151174
rect 257514 150854 258134 150938
rect 257514 150618 257546 150854
rect 257782 150618 257866 150854
rect 258102 150618 258134 150854
rect 257514 115174 258134 150618
rect 257514 114938 257546 115174
rect 257782 114938 257866 115174
rect 258102 114938 258134 115174
rect 257514 114854 258134 114938
rect 257514 114618 257546 114854
rect 257782 114618 257866 114854
rect 258102 114618 258134 114854
rect 257514 79174 258134 114618
rect 257514 78938 257546 79174
rect 257782 78938 257866 79174
rect 258102 78938 258134 79174
rect 257514 78854 258134 78938
rect 257514 78618 257546 78854
rect 257782 78618 257866 78854
rect 258102 78618 258134 78854
rect 257514 43174 258134 78618
rect 257514 42938 257546 43174
rect 257782 42938 257866 43174
rect 258102 42938 258134 43174
rect 257514 42854 258134 42938
rect 257514 42618 257546 42854
rect 257782 42618 257866 42854
rect 258102 42618 258134 42854
rect 257514 7174 258134 42618
rect 257514 6938 257546 7174
rect 257782 6938 257866 7174
rect 258102 6938 258134 7174
rect 257514 6854 258134 6938
rect 257514 6618 257546 6854
rect 257782 6618 257866 6854
rect 258102 6618 258134 6854
rect 257514 -2266 258134 6618
rect 257514 -2502 257546 -2266
rect 257782 -2502 257866 -2266
rect 258102 -2502 258134 -2266
rect 257514 -2586 258134 -2502
rect 257514 -2822 257546 -2586
rect 257782 -2822 257866 -2586
rect 258102 -2822 258134 -2586
rect 257514 -3814 258134 -2822
rect 261234 190894 261854 198800
rect 261234 190658 261266 190894
rect 261502 190658 261586 190894
rect 261822 190658 261854 190894
rect 261234 190574 261854 190658
rect 261234 190338 261266 190574
rect 261502 190338 261586 190574
rect 261822 190338 261854 190574
rect 261234 154894 261854 190338
rect 261234 154658 261266 154894
rect 261502 154658 261586 154894
rect 261822 154658 261854 154894
rect 261234 154574 261854 154658
rect 261234 154338 261266 154574
rect 261502 154338 261586 154574
rect 261822 154338 261854 154574
rect 261234 118894 261854 154338
rect 261234 118658 261266 118894
rect 261502 118658 261586 118894
rect 261822 118658 261854 118894
rect 261234 118574 261854 118658
rect 261234 118338 261266 118574
rect 261502 118338 261586 118574
rect 261822 118338 261854 118574
rect 261234 82894 261854 118338
rect 261234 82658 261266 82894
rect 261502 82658 261586 82894
rect 261822 82658 261854 82894
rect 261234 82574 261854 82658
rect 261234 82338 261266 82574
rect 261502 82338 261586 82574
rect 261822 82338 261854 82574
rect 261234 46894 261854 82338
rect 261234 46658 261266 46894
rect 261502 46658 261586 46894
rect 261822 46658 261854 46894
rect 261234 46574 261854 46658
rect 261234 46338 261266 46574
rect 261502 46338 261586 46574
rect 261822 46338 261854 46574
rect 261234 10894 261854 46338
rect 261234 10658 261266 10894
rect 261502 10658 261586 10894
rect 261822 10658 261854 10894
rect 261234 10574 261854 10658
rect 261234 10338 261266 10574
rect 261502 10338 261586 10574
rect 261822 10338 261854 10574
rect 261234 -4186 261854 10338
rect 261234 -4422 261266 -4186
rect 261502 -4422 261586 -4186
rect 261822 -4422 261854 -4186
rect 261234 -4506 261854 -4422
rect 261234 -4742 261266 -4506
rect 261502 -4742 261586 -4506
rect 261822 -4742 261854 -4506
rect 261234 -5734 261854 -4742
rect 264954 194614 265574 198800
rect 264954 194378 264986 194614
rect 265222 194378 265306 194614
rect 265542 194378 265574 194614
rect 264954 194294 265574 194378
rect 264954 194058 264986 194294
rect 265222 194058 265306 194294
rect 265542 194058 265574 194294
rect 264954 158614 265574 194058
rect 264954 158378 264986 158614
rect 265222 158378 265306 158614
rect 265542 158378 265574 158614
rect 264954 158294 265574 158378
rect 264954 158058 264986 158294
rect 265222 158058 265306 158294
rect 265542 158058 265574 158294
rect 264954 122614 265574 158058
rect 264954 122378 264986 122614
rect 265222 122378 265306 122614
rect 265542 122378 265574 122614
rect 264954 122294 265574 122378
rect 264954 122058 264986 122294
rect 265222 122058 265306 122294
rect 265542 122058 265574 122294
rect 264954 86614 265574 122058
rect 264954 86378 264986 86614
rect 265222 86378 265306 86614
rect 265542 86378 265574 86614
rect 264954 86294 265574 86378
rect 264954 86058 264986 86294
rect 265222 86058 265306 86294
rect 265542 86058 265574 86294
rect 264954 50614 265574 86058
rect 264954 50378 264986 50614
rect 265222 50378 265306 50614
rect 265542 50378 265574 50614
rect 264954 50294 265574 50378
rect 264954 50058 264986 50294
rect 265222 50058 265306 50294
rect 265542 50058 265574 50294
rect 264954 14614 265574 50058
rect 264954 14378 264986 14614
rect 265222 14378 265306 14614
rect 265542 14378 265574 14614
rect 264954 14294 265574 14378
rect 264954 14058 264986 14294
rect 265222 14058 265306 14294
rect 265542 14058 265574 14294
rect 246954 -7302 246986 -7066
rect 247222 -7302 247306 -7066
rect 247542 -7302 247574 -7066
rect 246954 -7386 247574 -7302
rect 246954 -7622 246986 -7386
rect 247222 -7622 247306 -7386
rect 247542 -7622 247574 -7386
rect 246954 -7654 247574 -7622
rect 264954 -6106 265574 14058
rect 271794 165454 272414 198800
rect 271794 165218 271826 165454
rect 272062 165218 272146 165454
rect 272382 165218 272414 165454
rect 271794 165134 272414 165218
rect 271794 164898 271826 165134
rect 272062 164898 272146 165134
rect 272382 164898 272414 165134
rect 271794 129454 272414 164898
rect 271794 129218 271826 129454
rect 272062 129218 272146 129454
rect 272382 129218 272414 129454
rect 271794 129134 272414 129218
rect 271794 128898 271826 129134
rect 272062 128898 272146 129134
rect 272382 128898 272414 129134
rect 271794 93454 272414 128898
rect 271794 93218 271826 93454
rect 272062 93218 272146 93454
rect 272382 93218 272414 93454
rect 271794 93134 272414 93218
rect 271794 92898 271826 93134
rect 272062 92898 272146 93134
rect 272382 92898 272414 93134
rect 271794 57454 272414 92898
rect 271794 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 272414 57454
rect 271794 57134 272414 57218
rect 271794 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 272414 57134
rect 271794 21454 272414 56898
rect 271794 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 272414 21454
rect 271794 21134 272414 21218
rect 271794 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 272414 21134
rect 271794 -1306 272414 20898
rect 271794 -1542 271826 -1306
rect 272062 -1542 272146 -1306
rect 272382 -1542 272414 -1306
rect 271794 -1626 272414 -1542
rect 271794 -1862 271826 -1626
rect 272062 -1862 272146 -1626
rect 272382 -1862 272414 -1626
rect 271794 -1894 272414 -1862
rect 275514 169174 276134 198800
rect 275514 168938 275546 169174
rect 275782 168938 275866 169174
rect 276102 168938 276134 169174
rect 275514 168854 276134 168938
rect 275514 168618 275546 168854
rect 275782 168618 275866 168854
rect 276102 168618 276134 168854
rect 275514 133174 276134 168618
rect 275514 132938 275546 133174
rect 275782 132938 275866 133174
rect 276102 132938 276134 133174
rect 275514 132854 276134 132938
rect 275514 132618 275546 132854
rect 275782 132618 275866 132854
rect 276102 132618 276134 132854
rect 275514 97174 276134 132618
rect 275514 96938 275546 97174
rect 275782 96938 275866 97174
rect 276102 96938 276134 97174
rect 275514 96854 276134 96938
rect 275514 96618 275546 96854
rect 275782 96618 275866 96854
rect 276102 96618 276134 96854
rect 275514 61174 276134 96618
rect 275514 60938 275546 61174
rect 275782 60938 275866 61174
rect 276102 60938 276134 61174
rect 275514 60854 276134 60938
rect 275514 60618 275546 60854
rect 275782 60618 275866 60854
rect 276102 60618 276134 60854
rect 275514 25174 276134 60618
rect 275514 24938 275546 25174
rect 275782 24938 275866 25174
rect 276102 24938 276134 25174
rect 275514 24854 276134 24938
rect 275514 24618 275546 24854
rect 275782 24618 275866 24854
rect 276102 24618 276134 24854
rect 275514 -3226 276134 24618
rect 275514 -3462 275546 -3226
rect 275782 -3462 275866 -3226
rect 276102 -3462 276134 -3226
rect 275514 -3546 276134 -3462
rect 275514 -3782 275546 -3546
rect 275782 -3782 275866 -3546
rect 276102 -3782 276134 -3546
rect 275514 -3814 276134 -3782
rect 279234 172894 279854 198800
rect 279234 172658 279266 172894
rect 279502 172658 279586 172894
rect 279822 172658 279854 172894
rect 279234 172574 279854 172658
rect 279234 172338 279266 172574
rect 279502 172338 279586 172574
rect 279822 172338 279854 172574
rect 279234 136894 279854 172338
rect 279234 136658 279266 136894
rect 279502 136658 279586 136894
rect 279822 136658 279854 136894
rect 279234 136574 279854 136658
rect 279234 136338 279266 136574
rect 279502 136338 279586 136574
rect 279822 136338 279854 136574
rect 279234 100894 279854 136338
rect 279234 100658 279266 100894
rect 279502 100658 279586 100894
rect 279822 100658 279854 100894
rect 279234 100574 279854 100658
rect 279234 100338 279266 100574
rect 279502 100338 279586 100574
rect 279822 100338 279854 100574
rect 279234 64894 279854 100338
rect 279234 64658 279266 64894
rect 279502 64658 279586 64894
rect 279822 64658 279854 64894
rect 279234 64574 279854 64658
rect 279234 64338 279266 64574
rect 279502 64338 279586 64574
rect 279822 64338 279854 64574
rect 279234 28894 279854 64338
rect 279234 28658 279266 28894
rect 279502 28658 279586 28894
rect 279822 28658 279854 28894
rect 279234 28574 279854 28658
rect 279234 28338 279266 28574
rect 279502 28338 279586 28574
rect 279822 28338 279854 28574
rect 279234 -5146 279854 28338
rect 279234 -5382 279266 -5146
rect 279502 -5382 279586 -5146
rect 279822 -5382 279854 -5146
rect 279234 -5466 279854 -5382
rect 279234 -5702 279266 -5466
rect 279502 -5702 279586 -5466
rect 279822 -5702 279854 -5466
rect 279234 -5734 279854 -5702
rect 282954 176614 283574 198800
rect 282954 176378 282986 176614
rect 283222 176378 283306 176614
rect 283542 176378 283574 176614
rect 282954 176294 283574 176378
rect 282954 176058 282986 176294
rect 283222 176058 283306 176294
rect 283542 176058 283574 176294
rect 282954 140614 283574 176058
rect 282954 140378 282986 140614
rect 283222 140378 283306 140614
rect 283542 140378 283574 140614
rect 282954 140294 283574 140378
rect 282954 140058 282986 140294
rect 283222 140058 283306 140294
rect 283542 140058 283574 140294
rect 282954 104614 283574 140058
rect 282954 104378 282986 104614
rect 283222 104378 283306 104614
rect 283542 104378 283574 104614
rect 282954 104294 283574 104378
rect 282954 104058 282986 104294
rect 283222 104058 283306 104294
rect 283542 104058 283574 104294
rect 282954 68614 283574 104058
rect 282954 68378 282986 68614
rect 283222 68378 283306 68614
rect 283542 68378 283574 68614
rect 282954 68294 283574 68378
rect 282954 68058 282986 68294
rect 283222 68058 283306 68294
rect 283542 68058 283574 68294
rect 282954 32614 283574 68058
rect 282954 32378 282986 32614
rect 283222 32378 283306 32614
rect 283542 32378 283574 32614
rect 282954 32294 283574 32378
rect 282954 32058 282986 32294
rect 283222 32058 283306 32294
rect 283542 32058 283574 32294
rect 264954 -6342 264986 -6106
rect 265222 -6342 265306 -6106
rect 265542 -6342 265574 -6106
rect 264954 -6426 265574 -6342
rect 264954 -6662 264986 -6426
rect 265222 -6662 265306 -6426
rect 265542 -6662 265574 -6426
rect 264954 -7654 265574 -6662
rect 282954 -7066 283574 32058
rect 289794 183454 290414 198800
rect 289794 183218 289826 183454
rect 290062 183218 290146 183454
rect 290382 183218 290414 183454
rect 289794 183134 290414 183218
rect 289794 182898 289826 183134
rect 290062 182898 290146 183134
rect 290382 182898 290414 183134
rect 289794 147454 290414 182898
rect 289794 147218 289826 147454
rect 290062 147218 290146 147454
rect 290382 147218 290414 147454
rect 289794 147134 290414 147218
rect 289794 146898 289826 147134
rect 290062 146898 290146 147134
rect 290382 146898 290414 147134
rect 289794 111454 290414 146898
rect 289794 111218 289826 111454
rect 290062 111218 290146 111454
rect 290382 111218 290414 111454
rect 289794 111134 290414 111218
rect 289794 110898 289826 111134
rect 290062 110898 290146 111134
rect 290382 110898 290414 111134
rect 289794 75454 290414 110898
rect 289794 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 290414 75454
rect 289794 75134 290414 75218
rect 289794 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 290414 75134
rect 289794 39454 290414 74898
rect 289794 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 290414 39454
rect 289794 39134 290414 39218
rect 289794 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 290414 39134
rect 289794 3454 290414 38898
rect 289794 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 290414 3454
rect 289794 3134 290414 3218
rect 289794 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 290414 3134
rect 289794 -346 290414 2898
rect 289794 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 290414 -346
rect 289794 -666 290414 -582
rect 289794 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 290414 -666
rect 289794 -1894 290414 -902
rect 293514 187174 294134 198800
rect 293514 186938 293546 187174
rect 293782 186938 293866 187174
rect 294102 186938 294134 187174
rect 293514 186854 294134 186938
rect 293514 186618 293546 186854
rect 293782 186618 293866 186854
rect 294102 186618 294134 186854
rect 293514 151174 294134 186618
rect 293514 150938 293546 151174
rect 293782 150938 293866 151174
rect 294102 150938 294134 151174
rect 293514 150854 294134 150938
rect 293514 150618 293546 150854
rect 293782 150618 293866 150854
rect 294102 150618 294134 150854
rect 293514 115174 294134 150618
rect 293514 114938 293546 115174
rect 293782 114938 293866 115174
rect 294102 114938 294134 115174
rect 293514 114854 294134 114938
rect 293514 114618 293546 114854
rect 293782 114618 293866 114854
rect 294102 114618 294134 114854
rect 293514 79174 294134 114618
rect 293514 78938 293546 79174
rect 293782 78938 293866 79174
rect 294102 78938 294134 79174
rect 293514 78854 294134 78938
rect 293514 78618 293546 78854
rect 293782 78618 293866 78854
rect 294102 78618 294134 78854
rect 293514 43174 294134 78618
rect 293514 42938 293546 43174
rect 293782 42938 293866 43174
rect 294102 42938 294134 43174
rect 293514 42854 294134 42938
rect 293514 42618 293546 42854
rect 293782 42618 293866 42854
rect 294102 42618 294134 42854
rect 293514 7174 294134 42618
rect 293514 6938 293546 7174
rect 293782 6938 293866 7174
rect 294102 6938 294134 7174
rect 293514 6854 294134 6938
rect 293514 6618 293546 6854
rect 293782 6618 293866 6854
rect 294102 6618 294134 6854
rect 293514 -2266 294134 6618
rect 293514 -2502 293546 -2266
rect 293782 -2502 293866 -2266
rect 294102 -2502 294134 -2266
rect 293514 -2586 294134 -2502
rect 293514 -2822 293546 -2586
rect 293782 -2822 293866 -2586
rect 294102 -2822 294134 -2586
rect 293514 -3814 294134 -2822
rect 297234 190894 297854 198800
rect 297234 190658 297266 190894
rect 297502 190658 297586 190894
rect 297822 190658 297854 190894
rect 297234 190574 297854 190658
rect 297234 190338 297266 190574
rect 297502 190338 297586 190574
rect 297822 190338 297854 190574
rect 297234 154894 297854 190338
rect 297234 154658 297266 154894
rect 297502 154658 297586 154894
rect 297822 154658 297854 154894
rect 297234 154574 297854 154658
rect 297234 154338 297266 154574
rect 297502 154338 297586 154574
rect 297822 154338 297854 154574
rect 297234 118894 297854 154338
rect 297234 118658 297266 118894
rect 297502 118658 297586 118894
rect 297822 118658 297854 118894
rect 297234 118574 297854 118658
rect 297234 118338 297266 118574
rect 297502 118338 297586 118574
rect 297822 118338 297854 118574
rect 297234 82894 297854 118338
rect 297234 82658 297266 82894
rect 297502 82658 297586 82894
rect 297822 82658 297854 82894
rect 297234 82574 297854 82658
rect 297234 82338 297266 82574
rect 297502 82338 297586 82574
rect 297822 82338 297854 82574
rect 297234 46894 297854 82338
rect 297234 46658 297266 46894
rect 297502 46658 297586 46894
rect 297822 46658 297854 46894
rect 297234 46574 297854 46658
rect 297234 46338 297266 46574
rect 297502 46338 297586 46574
rect 297822 46338 297854 46574
rect 297234 10894 297854 46338
rect 297234 10658 297266 10894
rect 297502 10658 297586 10894
rect 297822 10658 297854 10894
rect 297234 10574 297854 10658
rect 297234 10338 297266 10574
rect 297502 10338 297586 10574
rect 297822 10338 297854 10574
rect 297234 -4186 297854 10338
rect 297234 -4422 297266 -4186
rect 297502 -4422 297586 -4186
rect 297822 -4422 297854 -4186
rect 297234 -4506 297854 -4422
rect 297234 -4742 297266 -4506
rect 297502 -4742 297586 -4506
rect 297822 -4742 297854 -4506
rect 297234 -5734 297854 -4742
rect 300954 194614 301574 198800
rect 300954 194378 300986 194614
rect 301222 194378 301306 194614
rect 301542 194378 301574 194614
rect 300954 194294 301574 194378
rect 300954 194058 300986 194294
rect 301222 194058 301306 194294
rect 301542 194058 301574 194294
rect 300954 158614 301574 194058
rect 300954 158378 300986 158614
rect 301222 158378 301306 158614
rect 301542 158378 301574 158614
rect 300954 158294 301574 158378
rect 300954 158058 300986 158294
rect 301222 158058 301306 158294
rect 301542 158058 301574 158294
rect 300954 122614 301574 158058
rect 300954 122378 300986 122614
rect 301222 122378 301306 122614
rect 301542 122378 301574 122614
rect 300954 122294 301574 122378
rect 300954 122058 300986 122294
rect 301222 122058 301306 122294
rect 301542 122058 301574 122294
rect 300954 86614 301574 122058
rect 300954 86378 300986 86614
rect 301222 86378 301306 86614
rect 301542 86378 301574 86614
rect 300954 86294 301574 86378
rect 300954 86058 300986 86294
rect 301222 86058 301306 86294
rect 301542 86058 301574 86294
rect 300954 50614 301574 86058
rect 300954 50378 300986 50614
rect 301222 50378 301306 50614
rect 301542 50378 301574 50614
rect 300954 50294 301574 50378
rect 300954 50058 300986 50294
rect 301222 50058 301306 50294
rect 301542 50058 301574 50294
rect 300954 14614 301574 50058
rect 300954 14378 300986 14614
rect 301222 14378 301306 14614
rect 301542 14378 301574 14614
rect 300954 14294 301574 14378
rect 300954 14058 300986 14294
rect 301222 14058 301306 14294
rect 301542 14058 301574 14294
rect 282954 -7302 282986 -7066
rect 283222 -7302 283306 -7066
rect 283542 -7302 283574 -7066
rect 282954 -7386 283574 -7302
rect 282954 -7622 282986 -7386
rect 283222 -7622 283306 -7386
rect 283542 -7622 283574 -7386
rect 282954 -7654 283574 -7622
rect 300954 -6106 301574 14058
rect 307794 165454 308414 198800
rect 307794 165218 307826 165454
rect 308062 165218 308146 165454
rect 308382 165218 308414 165454
rect 307794 165134 308414 165218
rect 307794 164898 307826 165134
rect 308062 164898 308146 165134
rect 308382 164898 308414 165134
rect 307794 129454 308414 164898
rect 307794 129218 307826 129454
rect 308062 129218 308146 129454
rect 308382 129218 308414 129454
rect 307794 129134 308414 129218
rect 307794 128898 307826 129134
rect 308062 128898 308146 129134
rect 308382 128898 308414 129134
rect 307794 93454 308414 128898
rect 307794 93218 307826 93454
rect 308062 93218 308146 93454
rect 308382 93218 308414 93454
rect 307794 93134 308414 93218
rect 307794 92898 307826 93134
rect 308062 92898 308146 93134
rect 308382 92898 308414 93134
rect 307794 57454 308414 92898
rect 307794 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 308414 57454
rect 307794 57134 308414 57218
rect 307794 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 308414 57134
rect 307794 21454 308414 56898
rect 307794 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 308414 21454
rect 307794 21134 308414 21218
rect 307794 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 308414 21134
rect 307794 -1306 308414 20898
rect 307794 -1542 307826 -1306
rect 308062 -1542 308146 -1306
rect 308382 -1542 308414 -1306
rect 307794 -1626 308414 -1542
rect 307794 -1862 307826 -1626
rect 308062 -1862 308146 -1626
rect 308382 -1862 308414 -1626
rect 307794 -1894 308414 -1862
rect 311514 169174 312134 198800
rect 311514 168938 311546 169174
rect 311782 168938 311866 169174
rect 312102 168938 312134 169174
rect 311514 168854 312134 168938
rect 311514 168618 311546 168854
rect 311782 168618 311866 168854
rect 312102 168618 312134 168854
rect 311514 133174 312134 168618
rect 311514 132938 311546 133174
rect 311782 132938 311866 133174
rect 312102 132938 312134 133174
rect 311514 132854 312134 132938
rect 311514 132618 311546 132854
rect 311782 132618 311866 132854
rect 312102 132618 312134 132854
rect 311514 97174 312134 132618
rect 311514 96938 311546 97174
rect 311782 96938 311866 97174
rect 312102 96938 312134 97174
rect 311514 96854 312134 96938
rect 311514 96618 311546 96854
rect 311782 96618 311866 96854
rect 312102 96618 312134 96854
rect 311514 61174 312134 96618
rect 311514 60938 311546 61174
rect 311782 60938 311866 61174
rect 312102 60938 312134 61174
rect 311514 60854 312134 60938
rect 311514 60618 311546 60854
rect 311782 60618 311866 60854
rect 312102 60618 312134 60854
rect 311514 25174 312134 60618
rect 311514 24938 311546 25174
rect 311782 24938 311866 25174
rect 312102 24938 312134 25174
rect 311514 24854 312134 24938
rect 311514 24618 311546 24854
rect 311782 24618 311866 24854
rect 312102 24618 312134 24854
rect 311514 -3226 312134 24618
rect 311514 -3462 311546 -3226
rect 311782 -3462 311866 -3226
rect 312102 -3462 312134 -3226
rect 311514 -3546 312134 -3462
rect 311514 -3782 311546 -3546
rect 311782 -3782 311866 -3546
rect 312102 -3782 312134 -3546
rect 311514 -3814 312134 -3782
rect 315234 172894 315854 198800
rect 315234 172658 315266 172894
rect 315502 172658 315586 172894
rect 315822 172658 315854 172894
rect 315234 172574 315854 172658
rect 315234 172338 315266 172574
rect 315502 172338 315586 172574
rect 315822 172338 315854 172574
rect 315234 136894 315854 172338
rect 315234 136658 315266 136894
rect 315502 136658 315586 136894
rect 315822 136658 315854 136894
rect 315234 136574 315854 136658
rect 315234 136338 315266 136574
rect 315502 136338 315586 136574
rect 315822 136338 315854 136574
rect 315234 100894 315854 136338
rect 315234 100658 315266 100894
rect 315502 100658 315586 100894
rect 315822 100658 315854 100894
rect 315234 100574 315854 100658
rect 315234 100338 315266 100574
rect 315502 100338 315586 100574
rect 315822 100338 315854 100574
rect 315234 64894 315854 100338
rect 315234 64658 315266 64894
rect 315502 64658 315586 64894
rect 315822 64658 315854 64894
rect 315234 64574 315854 64658
rect 315234 64338 315266 64574
rect 315502 64338 315586 64574
rect 315822 64338 315854 64574
rect 315234 28894 315854 64338
rect 315234 28658 315266 28894
rect 315502 28658 315586 28894
rect 315822 28658 315854 28894
rect 315234 28574 315854 28658
rect 315234 28338 315266 28574
rect 315502 28338 315586 28574
rect 315822 28338 315854 28574
rect 315234 -5146 315854 28338
rect 315234 -5382 315266 -5146
rect 315502 -5382 315586 -5146
rect 315822 -5382 315854 -5146
rect 315234 -5466 315854 -5382
rect 315234 -5702 315266 -5466
rect 315502 -5702 315586 -5466
rect 315822 -5702 315854 -5466
rect 315234 -5734 315854 -5702
rect 318954 176614 319574 198800
rect 318954 176378 318986 176614
rect 319222 176378 319306 176614
rect 319542 176378 319574 176614
rect 318954 176294 319574 176378
rect 318954 176058 318986 176294
rect 319222 176058 319306 176294
rect 319542 176058 319574 176294
rect 318954 140614 319574 176058
rect 318954 140378 318986 140614
rect 319222 140378 319306 140614
rect 319542 140378 319574 140614
rect 318954 140294 319574 140378
rect 318954 140058 318986 140294
rect 319222 140058 319306 140294
rect 319542 140058 319574 140294
rect 318954 104614 319574 140058
rect 318954 104378 318986 104614
rect 319222 104378 319306 104614
rect 319542 104378 319574 104614
rect 318954 104294 319574 104378
rect 318954 104058 318986 104294
rect 319222 104058 319306 104294
rect 319542 104058 319574 104294
rect 318954 68614 319574 104058
rect 318954 68378 318986 68614
rect 319222 68378 319306 68614
rect 319542 68378 319574 68614
rect 318954 68294 319574 68378
rect 318954 68058 318986 68294
rect 319222 68058 319306 68294
rect 319542 68058 319574 68294
rect 318954 32614 319574 68058
rect 318954 32378 318986 32614
rect 319222 32378 319306 32614
rect 319542 32378 319574 32614
rect 318954 32294 319574 32378
rect 318954 32058 318986 32294
rect 319222 32058 319306 32294
rect 319542 32058 319574 32294
rect 300954 -6342 300986 -6106
rect 301222 -6342 301306 -6106
rect 301542 -6342 301574 -6106
rect 300954 -6426 301574 -6342
rect 300954 -6662 300986 -6426
rect 301222 -6662 301306 -6426
rect 301542 -6662 301574 -6426
rect 300954 -7654 301574 -6662
rect 318954 -7066 319574 32058
rect 325794 183454 326414 198800
rect 325794 183218 325826 183454
rect 326062 183218 326146 183454
rect 326382 183218 326414 183454
rect 325794 183134 326414 183218
rect 325794 182898 325826 183134
rect 326062 182898 326146 183134
rect 326382 182898 326414 183134
rect 325794 147454 326414 182898
rect 325794 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 326414 147454
rect 325794 147134 326414 147218
rect 325794 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 326414 147134
rect 325794 111454 326414 146898
rect 325794 111218 325826 111454
rect 326062 111218 326146 111454
rect 326382 111218 326414 111454
rect 325794 111134 326414 111218
rect 325794 110898 325826 111134
rect 326062 110898 326146 111134
rect 326382 110898 326414 111134
rect 325794 75454 326414 110898
rect 325794 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 326414 75454
rect 325794 75134 326414 75218
rect 325794 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 326414 75134
rect 325794 39454 326414 74898
rect 325794 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 326414 39454
rect 325794 39134 326414 39218
rect 325794 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 326414 39134
rect 325794 3454 326414 38898
rect 325794 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 326414 3454
rect 325794 3134 326414 3218
rect 325794 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 326414 3134
rect 325794 -346 326414 2898
rect 325794 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 326414 -346
rect 325794 -666 326414 -582
rect 325794 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 326414 -666
rect 325794 -1894 326414 -902
rect 329514 187174 330134 198800
rect 329514 186938 329546 187174
rect 329782 186938 329866 187174
rect 330102 186938 330134 187174
rect 329514 186854 330134 186938
rect 329514 186618 329546 186854
rect 329782 186618 329866 186854
rect 330102 186618 330134 186854
rect 329514 151174 330134 186618
rect 329514 150938 329546 151174
rect 329782 150938 329866 151174
rect 330102 150938 330134 151174
rect 329514 150854 330134 150938
rect 329514 150618 329546 150854
rect 329782 150618 329866 150854
rect 330102 150618 330134 150854
rect 329514 115174 330134 150618
rect 329514 114938 329546 115174
rect 329782 114938 329866 115174
rect 330102 114938 330134 115174
rect 329514 114854 330134 114938
rect 329514 114618 329546 114854
rect 329782 114618 329866 114854
rect 330102 114618 330134 114854
rect 329514 79174 330134 114618
rect 329514 78938 329546 79174
rect 329782 78938 329866 79174
rect 330102 78938 330134 79174
rect 329514 78854 330134 78938
rect 329514 78618 329546 78854
rect 329782 78618 329866 78854
rect 330102 78618 330134 78854
rect 329514 43174 330134 78618
rect 329514 42938 329546 43174
rect 329782 42938 329866 43174
rect 330102 42938 330134 43174
rect 329514 42854 330134 42938
rect 329514 42618 329546 42854
rect 329782 42618 329866 42854
rect 330102 42618 330134 42854
rect 329514 7174 330134 42618
rect 329514 6938 329546 7174
rect 329782 6938 329866 7174
rect 330102 6938 330134 7174
rect 329514 6854 330134 6938
rect 329514 6618 329546 6854
rect 329782 6618 329866 6854
rect 330102 6618 330134 6854
rect 329514 -2266 330134 6618
rect 329514 -2502 329546 -2266
rect 329782 -2502 329866 -2266
rect 330102 -2502 330134 -2266
rect 329514 -2586 330134 -2502
rect 329514 -2822 329546 -2586
rect 329782 -2822 329866 -2586
rect 330102 -2822 330134 -2586
rect 329514 -3814 330134 -2822
rect 333234 190894 333854 198800
rect 333234 190658 333266 190894
rect 333502 190658 333586 190894
rect 333822 190658 333854 190894
rect 333234 190574 333854 190658
rect 333234 190338 333266 190574
rect 333502 190338 333586 190574
rect 333822 190338 333854 190574
rect 333234 154894 333854 190338
rect 333234 154658 333266 154894
rect 333502 154658 333586 154894
rect 333822 154658 333854 154894
rect 333234 154574 333854 154658
rect 333234 154338 333266 154574
rect 333502 154338 333586 154574
rect 333822 154338 333854 154574
rect 333234 118894 333854 154338
rect 333234 118658 333266 118894
rect 333502 118658 333586 118894
rect 333822 118658 333854 118894
rect 333234 118574 333854 118658
rect 333234 118338 333266 118574
rect 333502 118338 333586 118574
rect 333822 118338 333854 118574
rect 333234 82894 333854 118338
rect 333234 82658 333266 82894
rect 333502 82658 333586 82894
rect 333822 82658 333854 82894
rect 333234 82574 333854 82658
rect 333234 82338 333266 82574
rect 333502 82338 333586 82574
rect 333822 82338 333854 82574
rect 333234 46894 333854 82338
rect 333234 46658 333266 46894
rect 333502 46658 333586 46894
rect 333822 46658 333854 46894
rect 333234 46574 333854 46658
rect 333234 46338 333266 46574
rect 333502 46338 333586 46574
rect 333822 46338 333854 46574
rect 333234 10894 333854 46338
rect 333234 10658 333266 10894
rect 333502 10658 333586 10894
rect 333822 10658 333854 10894
rect 333234 10574 333854 10658
rect 333234 10338 333266 10574
rect 333502 10338 333586 10574
rect 333822 10338 333854 10574
rect 333234 -4186 333854 10338
rect 333234 -4422 333266 -4186
rect 333502 -4422 333586 -4186
rect 333822 -4422 333854 -4186
rect 333234 -4506 333854 -4422
rect 333234 -4742 333266 -4506
rect 333502 -4742 333586 -4506
rect 333822 -4742 333854 -4506
rect 333234 -5734 333854 -4742
rect 336954 194614 337574 198800
rect 336954 194378 336986 194614
rect 337222 194378 337306 194614
rect 337542 194378 337574 194614
rect 336954 194294 337574 194378
rect 336954 194058 336986 194294
rect 337222 194058 337306 194294
rect 337542 194058 337574 194294
rect 336954 158614 337574 194058
rect 336954 158378 336986 158614
rect 337222 158378 337306 158614
rect 337542 158378 337574 158614
rect 336954 158294 337574 158378
rect 336954 158058 336986 158294
rect 337222 158058 337306 158294
rect 337542 158058 337574 158294
rect 336954 122614 337574 158058
rect 336954 122378 336986 122614
rect 337222 122378 337306 122614
rect 337542 122378 337574 122614
rect 336954 122294 337574 122378
rect 336954 122058 336986 122294
rect 337222 122058 337306 122294
rect 337542 122058 337574 122294
rect 336954 86614 337574 122058
rect 336954 86378 336986 86614
rect 337222 86378 337306 86614
rect 337542 86378 337574 86614
rect 336954 86294 337574 86378
rect 336954 86058 336986 86294
rect 337222 86058 337306 86294
rect 337542 86058 337574 86294
rect 336954 50614 337574 86058
rect 336954 50378 336986 50614
rect 337222 50378 337306 50614
rect 337542 50378 337574 50614
rect 336954 50294 337574 50378
rect 336954 50058 336986 50294
rect 337222 50058 337306 50294
rect 337542 50058 337574 50294
rect 336954 14614 337574 50058
rect 336954 14378 336986 14614
rect 337222 14378 337306 14614
rect 337542 14378 337574 14614
rect 336954 14294 337574 14378
rect 336954 14058 336986 14294
rect 337222 14058 337306 14294
rect 337542 14058 337574 14294
rect 318954 -7302 318986 -7066
rect 319222 -7302 319306 -7066
rect 319542 -7302 319574 -7066
rect 318954 -7386 319574 -7302
rect 318954 -7622 318986 -7386
rect 319222 -7622 319306 -7386
rect 319542 -7622 319574 -7386
rect 318954 -7654 319574 -7622
rect 336954 -6106 337574 14058
rect 343794 165454 344414 198800
rect 343794 165218 343826 165454
rect 344062 165218 344146 165454
rect 344382 165218 344414 165454
rect 343794 165134 344414 165218
rect 343794 164898 343826 165134
rect 344062 164898 344146 165134
rect 344382 164898 344414 165134
rect 343794 129454 344414 164898
rect 343794 129218 343826 129454
rect 344062 129218 344146 129454
rect 344382 129218 344414 129454
rect 343794 129134 344414 129218
rect 343794 128898 343826 129134
rect 344062 128898 344146 129134
rect 344382 128898 344414 129134
rect 343794 93454 344414 128898
rect 343794 93218 343826 93454
rect 344062 93218 344146 93454
rect 344382 93218 344414 93454
rect 343794 93134 344414 93218
rect 343794 92898 343826 93134
rect 344062 92898 344146 93134
rect 344382 92898 344414 93134
rect 343794 57454 344414 92898
rect 343794 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 344414 57454
rect 343794 57134 344414 57218
rect 343794 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 344414 57134
rect 343794 21454 344414 56898
rect 343794 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 344414 21454
rect 343794 21134 344414 21218
rect 343794 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 344414 21134
rect 343794 -1306 344414 20898
rect 343794 -1542 343826 -1306
rect 344062 -1542 344146 -1306
rect 344382 -1542 344414 -1306
rect 343794 -1626 344414 -1542
rect 343794 -1862 343826 -1626
rect 344062 -1862 344146 -1626
rect 344382 -1862 344414 -1626
rect 343794 -1894 344414 -1862
rect 347514 169174 348134 198800
rect 347514 168938 347546 169174
rect 347782 168938 347866 169174
rect 348102 168938 348134 169174
rect 347514 168854 348134 168938
rect 347514 168618 347546 168854
rect 347782 168618 347866 168854
rect 348102 168618 348134 168854
rect 347514 133174 348134 168618
rect 347514 132938 347546 133174
rect 347782 132938 347866 133174
rect 348102 132938 348134 133174
rect 347514 132854 348134 132938
rect 347514 132618 347546 132854
rect 347782 132618 347866 132854
rect 348102 132618 348134 132854
rect 347514 97174 348134 132618
rect 347514 96938 347546 97174
rect 347782 96938 347866 97174
rect 348102 96938 348134 97174
rect 347514 96854 348134 96938
rect 347514 96618 347546 96854
rect 347782 96618 347866 96854
rect 348102 96618 348134 96854
rect 347514 61174 348134 96618
rect 347514 60938 347546 61174
rect 347782 60938 347866 61174
rect 348102 60938 348134 61174
rect 347514 60854 348134 60938
rect 347514 60618 347546 60854
rect 347782 60618 347866 60854
rect 348102 60618 348134 60854
rect 347514 25174 348134 60618
rect 347514 24938 347546 25174
rect 347782 24938 347866 25174
rect 348102 24938 348134 25174
rect 347514 24854 348134 24938
rect 347514 24618 347546 24854
rect 347782 24618 347866 24854
rect 348102 24618 348134 24854
rect 347514 -3226 348134 24618
rect 347514 -3462 347546 -3226
rect 347782 -3462 347866 -3226
rect 348102 -3462 348134 -3226
rect 347514 -3546 348134 -3462
rect 347514 -3782 347546 -3546
rect 347782 -3782 347866 -3546
rect 348102 -3782 348134 -3546
rect 347514 -3814 348134 -3782
rect 351234 172894 351854 198800
rect 351234 172658 351266 172894
rect 351502 172658 351586 172894
rect 351822 172658 351854 172894
rect 351234 172574 351854 172658
rect 351234 172338 351266 172574
rect 351502 172338 351586 172574
rect 351822 172338 351854 172574
rect 351234 136894 351854 172338
rect 351234 136658 351266 136894
rect 351502 136658 351586 136894
rect 351822 136658 351854 136894
rect 351234 136574 351854 136658
rect 351234 136338 351266 136574
rect 351502 136338 351586 136574
rect 351822 136338 351854 136574
rect 351234 100894 351854 136338
rect 351234 100658 351266 100894
rect 351502 100658 351586 100894
rect 351822 100658 351854 100894
rect 351234 100574 351854 100658
rect 351234 100338 351266 100574
rect 351502 100338 351586 100574
rect 351822 100338 351854 100574
rect 351234 64894 351854 100338
rect 351234 64658 351266 64894
rect 351502 64658 351586 64894
rect 351822 64658 351854 64894
rect 351234 64574 351854 64658
rect 351234 64338 351266 64574
rect 351502 64338 351586 64574
rect 351822 64338 351854 64574
rect 351234 28894 351854 64338
rect 351234 28658 351266 28894
rect 351502 28658 351586 28894
rect 351822 28658 351854 28894
rect 351234 28574 351854 28658
rect 351234 28338 351266 28574
rect 351502 28338 351586 28574
rect 351822 28338 351854 28574
rect 351234 -5146 351854 28338
rect 351234 -5382 351266 -5146
rect 351502 -5382 351586 -5146
rect 351822 -5382 351854 -5146
rect 351234 -5466 351854 -5382
rect 351234 -5702 351266 -5466
rect 351502 -5702 351586 -5466
rect 351822 -5702 351854 -5466
rect 351234 -5734 351854 -5702
rect 354954 176614 355574 198800
rect 354954 176378 354986 176614
rect 355222 176378 355306 176614
rect 355542 176378 355574 176614
rect 354954 176294 355574 176378
rect 354954 176058 354986 176294
rect 355222 176058 355306 176294
rect 355542 176058 355574 176294
rect 354954 140614 355574 176058
rect 354954 140378 354986 140614
rect 355222 140378 355306 140614
rect 355542 140378 355574 140614
rect 354954 140294 355574 140378
rect 354954 140058 354986 140294
rect 355222 140058 355306 140294
rect 355542 140058 355574 140294
rect 354954 104614 355574 140058
rect 354954 104378 354986 104614
rect 355222 104378 355306 104614
rect 355542 104378 355574 104614
rect 354954 104294 355574 104378
rect 354954 104058 354986 104294
rect 355222 104058 355306 104294
rect 355542 104058 355574 104294
rect 354954 68614 355574 104058
rect 354954 68378 354986 68614
rect 355222 68378 355306 68614
rect 355542 68378 355574 68614
rect 354954 68294 355574 68378
rect 354954 68058 354986 68294
rect 355222 68058 355306 68294
rect 355542 68058 355574 68294
rect 354954 32614 355574 68058
rect 354954 32378 354986 32614
rect 355222 32378 355306 32614
rect 355542 32378 355574 32614
rect 354954 32294 355574 32378
rect 354954 32058 354986 32294
rect 355222 32058 355306 32294
rect 355542 32058 355574 32294
rect 336954 -6342 336986 -6106
rect 337222 -6342 337306 -6106
rect 337542 -6342 337574 -6106
rect 336954 -6426 337574 -6342
rect 336954 -6662 336986 -6426
rect 337222 -6662 337306 -6426
rect 337542 -6662 337574 -6426
rect 336954 -7654 337574 -6662
rect 354954 -7066 355574 32058
rect 361794 183454 362414 198800
rect 361794 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 362414 183454
rect 361794 183134 362414 183218
rect 361794 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 362414 183134
rect 361794 147454 362414 182898
rect 361794 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 362414 147454
rect 361794 147134 362414 147218
rect 361794 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 362414 147134
rect 361794 111454 362414 146898
rect 361794 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 362414 111454
rect 361794 111134 362414 111218
rect 361794 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 362414 111134
rect 361794 75454 362414 110898
rect 361794 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 362414 75454
rect 361794 75134 362414 75218
rect 361794 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 362414 75134
rect 361794 39454 362414 74898
rect 361794 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 362414 39454
rect 361794 39134 362414 39218
rect 361794 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 362414 39134
rect 361794 3454 362414 38898
rect 361794 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 362414 3454
rect 361794 3134 362414 3218
rect 361794 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 362414 3134
rect 361794 -346 362414 2898
rect 361794 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 362414 -346
rect 361794 -666 362414 -582
rect 361794 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 362414 -666
rect 361794 -1894 362414 -902
rect 365514 187174 366134 198800
rect 365514 186938 365546 187174
rect 365782 186938 365866 187174
rect 366102 186938 366134 187174
rect 365514 186854 366134 186938
rect 365514 186618 365546 186854
rect 365782 186618 365866 186854
rect 366102 186618 366134 186854
rect 365514 151174 366134 186618
rect 365514 150938 365546 151174
rect 365782 150938 365866 151174
rect 366102 150938 366134 151174
rect 365514 150854 366134 150938
rect 365514 150618 365546 150854
rect 365782 150618 365866 150854
rect 366102 150618 366134 150854
rect 365514 115174 366134 150618
rect 365514 114938 365546 115174
rect 365782 114938 365866 115174
rect 366102 114938 366134 115174
rect 365514 114854 366134 114938
rect 365514 114618 365546 114854
rect 365782 114618 365866 114854
rect 366102 114618 366134 114854
rect 365514 79174 366134 114618
rect 365514 78938 365546 79174
rect 365782 78938 365866 79174
rect 366102 78938 366134 79174
rect 365514 78854 366134 78938
rect 365514 78618 365546 78854
rect 365782 78618 365866 78854
rect 366102 78618 366134 78854
rect 365514 43174 366134 78618
rect 365514 42938 365546 43174
rect 365782 42938 365866 43174
rect 366102 42938 366134 43174
rect 365514 42854 366134 42938
rect 365514 42618 365546 42854
rect 365782 42618 365866 42854
rect 366102 42618 366134 42854
rect 365514 7174 366134 42618
rect 365514 6938 365546 7174
rect 365782 6938 365866 7174
rect 366102 6938 366134 7174
rect 365514 6854 366134 6938
rect 365514 6618 365546 6854
rect 365782 6618 365866 6854
rect 366102 6618 366134 6854
rect 365514 -2266 366134 6618
rect 365514 -2502 365546 -2266
rect 365782 -2502 365866 -2266
rect 366102 -2502 366134 -2266
rect 365514 -2586 366134 -2502
rect 365514 -2822 365546 -2586
rect 365782 -2822 365866 -2586
rect 366102 -2822 366134 -2586
rect 365514 -3814 366134 -2822
rect 369234 190894 369854 198800
rect 369234 190658 369266 190894
rect 369502 190658 369586 190894
rect 369822 190658 369854 190894
rect 369234 190574 369854 190658
rect 369234 190338 369266 190574
rect 369502 190338 369586 190574
rect 369822 190338 369854 190574
rect 369234 154894 369854 190338
rect 369234 154658 369266 154894
rect 369502 154658 369586 154894
rect 369822 154658 369854 154894
rect 369234 154574 369854 154658
rect 369234 154338 369266 154574
rect 369502 154338 369586 154574
rect 369822 154338 369854 154574
rect 369234 118894 369854 154338
rect 369234 118658 369266 118894
rect 369502 118658 369586 118894
rect 369822 118658 369854 118894
rect 369234 118574 369854 118658
rect 369234 118338 369266 118574
rect 369502 118338 369586 118574
rect 369822 118338 369854 118574
rect 369234 82894 369854 118338
rect 369234 82658 369266 82894
rect 369502 82658 369586 82894
rect 369822 82658 369854 82894
rect 369234 82574 369854 82658
rect 369234 82338 369266 82574
rect 369502 82338 369586 82574
rect 369822 82338 369854 82574
rect 369234 46894 369854 82338
rect 369234 46658 369266 46894
rect 369502 46658 369586 46894
rect 369822 46658 369854 46894
rect 369234 46574 369854 46658
rect 369234 46338 369266 46574
rect 369502 46338 369586 46574
rect 369822 46338 369854 46574
rect 369234 10894 369854 46338
rect 369234 10658 369266 10894
rect 369502 10658 369586 10894
rect 369822 10658 369854 10894
rect 369234 10574 369854 10658
rect 369234 10338 369266 10574
rect 369502 10338 369586 10574
rect 369822 10338 369854 10574
rect 369234 -4186 369854 10338
rect 369234 -4422 369266 -4186
rect 369502 -4422 369586 -4186
rect 369822 -4422 369854 -4186
rect 369234 -4506 369854 -4422
rect 369234 -4742 369266 -4506
rect 369502 -4742 369586 -4506
rect 369822 -4742 369854 -4506
rect 369234 -5734 369854 -4742
rect 372954 194614 373574 198800
rect 372954 194378 372986 194614
rect 373222 194378 373306 194614
rect 373542 194378 373574 194614
rect 372954 194294 373574 194378
rect 372954 194058 372986 194294
rect 373222 194058 373306 194294
rect 373542 194058 373574 194294
rect 372954 158614 373574 194058
rect 372954 158378 372986 158614
rect 373222 158378 373306 158614
rect 373542 158378 373574 158614
rect 372954 158294 373574 158378
rect 372954 158058 372986 158294
rect 373222 158058 373306 158294
rect 373542 158058 373574 158294
rect 372954 122614 373574 158058
rect 372954 122378 372986 122614
rect 373222 122378 373306 122614
rect 373542 122378 373574 122614
rect 372954 122294 373574 122378
rect 372954 122058 372986 122294
rect 373222 122058 373306 122294
rect 373542 122058 373574 122294
rect 372954 86614 373574 122058
rect 372954 86378 372986 86614
rect 373222 86378 373306 86614
rect 373542 86378 373574 86614
rect 372954 86294 373574 86378
rect 372954 86058 372986 86294
rect 373222 86058 373306 86294
rect 373542 86058 373574 86294
rect 372954 50614 373574 86058
rect 372954 50378 372986 50614
rect 373222 50378 373306 50614
rect 373542 50378 373574 50614
rect 372954 50294 373574 50378
rect 372954 50058 372986 50294
rect 373222 50058 373306 50294
rect 373542 50058 373574 50294
rect 372954 14614 373574 50058
rect 372954 14378 372986 14614
rect 373222 14378 373306 14614
rect 373542 14378 373574 14614
rect 372954 14294 373574 14378
rect 372954 14058 372986 14294
rect 373222 14058 373306 14294
rect 373542 14058 373574 14294
rect 354954 -7302 354986 -7066
rect 355222 -7302 355306 -7066
rect 355542 -7302 355574 -7066
rect 354954 -7386 355574 -7302
rect 354954 -7622 354986 -7386
rect 355222 -7622 355306 -7386
rect 355542 -7622 355574 -7386
rect 354954 -7654 355574 -7622
rect 372954 -6106 373574 14058
rect 379794 165454 380414 198800
rect 379794 165218 379826 165454
rect 380062 165218 380146 165454
rect 380382 165218 380414 165454
rect 379794 165134 380414 165218
rect 379794 164898 379826 165134
rect 380062 164898 380146 165134
rect 380382 164898 380414 165134
rect 379794 129454 380414 164898
rect 379794 129218 379826 129454
rect 380062 129218 380146 129454
rect 380382 129218 380414 129454
rect 379794 129134 380414 129218
rect 379794 128898 379826 129134
rect 380062 128898 380146 129134
rect 380382 128898 380414 129134
rect 379794 93454 380414 128898
rect 379794 93218 379826 93454
rect 380062 93218 380146 93454
rect 380382 93218 380414 93454
rect 379794 93134 380414 93218
rect 379794 92898 379826 93134
rect 380062 92898 380146 93134
rect 380382 92898 380414 93134
rect 379794 57454 380414 92898
rect 379794 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 380414 57454
rect 379794 57134 380414 57218
rect 379794 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 380414 57134
rect 379794 21454 380414 56898
rect 379794 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 380414 21454
rect 379794 21134 380414 21218
rect 379794 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 380414 21134
rect 379794 -1306 380414 20898
rect 379794 -1542 379826 -1306
rect 380062 -1542 380146 -1306
rect 380382 -1542 380414 -1306
rect 379794 -1626 380414 -1542
rect 379794 -1862 379826 -1626
rect 380062 -1862 380146 -1626
rect 380382 -1862 380414 -1626
rect 379794 -1894 380414 -1862
rect 383514 169174 384134 198800
rect 383514 168938 383546 169174
rect 383782 168938 383866 169174
rect 384102 168938 384134 169174
rect 383514 168854 384134 168938
rect 383514 168618 383546 168854
rect 383782 168618 383866 168854
rect 384102 168618 384134 168854
rect 383514 133174 384134 168618
rect 383514 132938 383546 133174
rect 383782 132938 383866 133174
rect 384102 132938 384134 133174
rect 383514 132854 384134 132938
rect 383514 132618 383546 132854
rect 383782 132618 383866 132854
rect 384102 132618 384134 132854
rect 383514 97174 384134 132618
rect 383514 96938 383546 97174
rect 383782 96938 383866 97174
rect 384102 96938 384134 97174
rect 383514 96854 384134 96938
rect 383514 96618 383546 96854
rect 383782 96618 383866 96854
rect 384102 96618 384134 96854
rect 383514 61174 384134 96618
rect 383514 60938 383546 61174
rect 383782 60938 383866 61174
rect 384102 60938 384134 61174
rect 383514 60854 384134 60938
rect 383514 60618 383546 60854
rect 383782 60618 383866 60854
rect 384102 60618 384134 60854
rect 383514 25174 384134 60618
rect 383514 24938 383546 25174
rect 383782 24938 383866 25174
rect 384102 24938 384134 25174
rect 383514 24854 384134 24938
rect 383514 24618 383546 24854
rect 383782 24618 383866 24854
rect 384102 24618 384134 24854
rect 383514 -3226 384134 24618
rect 383514 -3462 383546 -3226
rect 383782 -3462 383866 -3226
rect 384102 -3462 384134 -3226
rect 383514 -3546 384134 -3462
rect 383514 -3782 383546 -3546
rect 383782 -3782 383866 -3546
rect 384102 -3782 384134 -3546
rect 383514 -3814 384134 -3782
rect 387234 172894 387854 198800
rect 387234 172658 387266 172894
rect 387502 172658 387586 172894
rect 387822 172658 387854 172894
rect 387234 172574 387854 172658
rect 387234 172338 387266 172574
rect 387502 172338 387586 172574
rect 387822 172338 387854 172574
rect 387234 136894 387854 172338
rect 387234 136658 387266 136894
rect 387502 136658 387586 136894
rect 387822 136658 387854 136894
rect 387234 136574 387854 136658
rect 387234 136338 387266 136574
rect 387502 136338 387586 136574
rect 387822 136338 387854 136574
rect 387234 100894 387854 136338
rect 387234 100658 387266 100894
rect 387502 100658 387586 100894
rect 387822 100658 387854 100894
rect 387234 100574 387854 100658
rect 387234 100338 387266 100574
rect 387502 100338 387586 100574
rect 387822 100338 387854 100574
rect 387234 64894 387854 100338
rect 387234 64658 387266 64894
rect 387502 64658 387586 64894
rect 387822 64658 387854 64894
rect 387234 64574 387854 64658
rect 387234 64338 387266 64574
rect 387502 64338 387586 64574
rect 387822 64338 387854 64574
rect 387234 28894 387854 64338
rect 387234 28658 387266 28894
rect 387502 28658 387586 28894
rect 387822 28658 387854 28894
rect 387234 28574 387854 28658
rect 387234 28338 387266 28574
rect 387502 28338 387586 28574
rect 387822 28338 387854 28574
rect 387234 -5146 387854 28338
rect 387234 -5382 387266 -5146
rect 387502 -5382 387586 -5146
rect 387822 -5382 387854 -5146
rect 387234 -5466 387854 -5382
rect 387234 -5702 387266 -5466
rect 387502 -5702 387586 -5466
rect 387822 -5702 387854 -5466
rect 387234 -5734 387854 -5702
rect 390954 176614 391574 198800
rect 390954 176378 390986 176614
rect 391222 176378 391306 176614
rect 391542 176378 391574 176614
rect 390954 176294 391574 176378
rect 390954 176058 390986 176294
rect 391222 176058 391306 176294
rect 391542 176058 391574 176294
rect 390954 140614 391574 176058
rect 390954 140378 390986 140614
rect 391222 140378 391306 140614
rect 391542 140378 391574 140614
rect 390954 140294 391574 140378
rect 390954 140058 390986 140294
rect 391222 140058 391306 140294
rect 391542 140058 391574 140294
rect 390954 104614 391574 140058
rect 390954 104378 390986 104614
rect 391222 104378 391306 104614
rect 391542 104378 391574 104614
rect 390954 104294 391574 104378
rect 390954 104058 390986 104294
rect 391222 104058 391306 104294
rect 391542 104058 391574 104294
rect 390954 68614 391574 104058
rect 390954 68378 390986 68614
rect 391222 68378 391306 68614
rect 391542 68378 391574 68614
rect 390954 68294 391574 68378
rect 390954 68058 390986 68294
rect 391222 68058 391306 68294
rect 391542 68058 391574 68294
rect 390954 32614 391574 68058
rect 390954 32378 390986 32614
rect 391222 32378 391306 32614
rect 391542 32378 391574 32614
rect 390954 32294 391574 32378
rect 390954 32058 390986 32294
rect 391222 32058 391306 32294
rect 391542 32058 391574 32294
rect 372954 -6342 372986 -6106
rect 373222 -6342 373306 -6106
rect 373542 -6342 373574 -6106
rect 372954 -6426 373574 -6342
rect 372954 -6662 372986 -6426
rect 373222 -6662 373306 -6426
rect 373542 -6662 373574 -6426
rect 372954 -7654 373574 -6662
rect 390954 -7066 391574 32058
rect 397794 183454 398414 198800
rect 397794 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 398414 183454
rect 397794 183134 398414 183218
rect 397794 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 398414 183134
rect 397794 147454 398414 182898
rect 397794 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 398414 147454
rect 397794 147134 398414 147218
rect 397794 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 398414 147134
rect 397794 111454 398414 146898
rect 397794 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 398414 111454
rect 397794 111134 398414 111218
rect 397794 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 398414 111134
rect 397794 75454 398414 110898
rect 397794 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 398414 75454
rect 397794 75134 398414 75218
rect 397794 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 398414 75134
rect 397794 39454 398414 74898
rect 397794 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 398414 39454
rect 397794 39134 398414 39218
rect 397794 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 398414 39134
rect 397794 3454 398414 38898
rect 397794 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 398414 3454
rect 397794 3134 398414 3218
rect 397794 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 398414 3134
rect 397794 -346 398414 2898
rect 397794 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 398414 -346
rect 397794 -666 398414 -582
rect 397794 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 398414 -666
rect 397794 -1894 398414 -902
rect 401514 187174 402134 198800
rect 401514 186938 401546 187174
rect 401782 186938 401866 187174
rect 402102 186938 402134 187174
rect 401514 186854 402134 186938
rect 401514 186618 401546 186854
rect 401782 186618 401866 186854
rect 402102 186618 402134 186854
rect 401514 151174 402134 186618
rect 401514 150938 401546 151174
rect 401782 150938 401866 151174
rect 402102 150938 402134 151174
rect 401514 150854 402134 150938
rect 401514 150618 401546 150854
rect 401782 150618 401866 150854
rect 402102 150618 402134 150854
rect 401514 115174 402134 150618
rect 401514 114938 401546 115174
rect 401782 114938 401866 115174
rect 402102 114938 402134 115174
rect 401514 114854 402134 114938
rect 401514 114618 401546 114854
rect 401782 114618 401866 114854
rect 402102 114618 402134 114854
rect 401514 79174 402134 114618
rect 401514 78938 401546 79174
rect 401782 78938 401866 79174
rect 402102 78938 402134 79174
rect 401514 78854 402134 78938
rect 401514 78618 401546 78854
rect 401782 78618 401866 78854
rect 402102 78618 402134 78854
rect 401514 43174 402134 78618
rect 401514 42938 401546 43174
rect 401782 42938 401866 43174
rect 402102 42938 402134 43174
rect 401514 42854 402134 42938
rect 401514 42618 401546 42854
rect 401782 42618 401866 42854
rect 402102 42618 402134 42854
rect 401514 7174 402134 42618
rect 401514 6938 401546 7174
rect 401782 6938 401866 7174
rect 402102 6938 402134 7174
rect 401514 6854 402134 6938
rect 401514 6618 401546 6854
rect 401782 6618 401866 6854
rect 402102 6618 402134 6854
rect 401514 -2266 402134 6618
rect 401514 -2502 401546 -2266
rect 401782 -2502 401866 -2266
rect 402102 -2502 402134 -2266
rect 401514 -2586 402134 -2502
rect 401514 -2822 401546 -2586
rect 401782 -2822 401866 -2586
rect 402102 -2822 402134 -2586
rect 401514 -3814 402134 -2822
rect 405234 190894 405854 198800
rect 405234 190658 405266 190894
rect 405502 190658 405586 190894
rect 405822 190658 405854 190894
rect 405234 190574 405854 190658
rect 405234 190338 405266 190574
rect 405502 190338 405586 190574
rect 405822 190338 405854 190574
rect 405234 154894 405854 190338
rect 405234 154658 405266 154894
rect 405502 154658 405586 154894
rect 405822 154658 405854 154894
rect 405234 154574 405854 154658
rect 405234 154338 405266 154574
rect 405502 154338 405586 154574
rect 405822 154338 405854 154574
rect 405234 118894 405854 154338
rect 405234 118658 405266 118894
rect 405502 118658 405586 118894
rect 405822 118658 405854 118894
rect 405234 118574 405854 118658
rect 405234 118338 405266 118574
rect 405502 118338 405586 118574
rect 405822 118338 405854 118574
rect 405234 82894 405854 118338
rect 405234 82658 405266 82894
rect 405502 82658 405586 82894
rect 405822 82658 405854 82894
rect 405234 82574 405854 82658
rect 405234 82338 405266 82574
rect 405502 82338 405586 82574
rect 405822 82338 405854 82574
rect 405234 46894 405854 82338
rect 405234 46658 405266 46894
rect 405502 46658 405586 46894
rect 405822 46658 405854 46894
rect 405234 46574 405854 46658
rect 405234 46338 405266 46574
rect 405502 46338 405586 46574
rect 405822 46338 405854 46574
rect 405234 10894 405854 46338
rect 405234 10658 405266 10894
rect 405502 10658 405586 10894
rect 405822 10658 405854 10894
rect 405234 10574 405854 10658
rect 405234 10338 405266 10574
rect 405502 10338 405586 10574
rect 405822 10338 405854 10574
rect 405234 -4186 405854 10338
rect 405234 -4422 405266 -4186
rect 405502 -4422 405586 -4186
rect 405822 -4422 405854 -4186
rect 405234 -4506 405854 -4422
rect 405234 -4742 405266 -4506
rect 405502 -4742 405586 -4506
rect 405822 -4742 405854 -4506
rect 405234 -5734 405854 -4742
rect 408954 194614 409574 198800
rect 408954 194378 408986 194614
rect 409222 194378 409306 194614
rect 409542 194378 409574 194614
rect 408954 194294 409574 194378
rect 408954 194058 408986 194294
rect 409222 194058 409306 194294
rect 409542 194058 409574 194294
rect 408954 158614 409574 194058
rect 408954 158378 408986 158614
rect 409222 158378 409306 158614
rect 409542 158378 409574 158614
rect 408954 158294 409574 158378
rect 408954 158058 408986 158294
rect 409222 158058 409306 158294
rect 409542 158058 409574 158294
rect 408954 122614 409574 158058
rect 408954 122378 408986 122614
rect 409222 122378 409306 122614
rect 409542 122378 409574 122614
rect 408954 122294 409574 122378
rect 408954 122058 408986 122294
rect 409222 122058 409306 122294
rect 409542 122058 409574 122294
rect 408954 86614 409574 122058
rect 408954 86378 408986 86614
rect 409222 86378 409306 86614
rect 409542 86378 409574 86614
rect 408954 86294 409574 86378
rect 408954 86058 408986 86294
rect 409222 86058 409306 86294
rect 409542 86058 409574 86294
rect 408954 50614 409574 86058
rect 408954 50378 408986 50614
rect 409222 50378 409306 50614
rect 409542 50378 409574 50614
rect 408954 50294 409574 50378
rect 408954 50058 408986 50294
rect 409222 50058 409306 50294
rect 409542 50058 409574 50294
rect 408954 14614 409574 50058
rect 408954 14378 408986 14614
rect 409222 14378 409306 14614
rect 409542 14378 409574 14614
rect 408954 14294 409574 14378
rect 408954 14058 408986 14294
rect 409222 14058 409306 14294
rect 409542 14058 409574 14294
rect 390954 -7302 390986 -7066
rect 391222 -7302 391306 -7066
rect 391542 -7302 391574 -7066
rect 390954 -7386 391574 -7302
rect 390954 -7622 390986 -7386
rect 391222 -7622 391306 -7386
rect 391542 -7622 391574 -7386
rect 390954 -7654 391574 -7622
rect 408954 -6106 409574 14058
rect 415794 165454 416414 198800
rect 415794 165218 415826 165454
rect 416062 165218 416146 165454
rect 416382 165218 416414 165454
rect 415794 165134 416414 165218
rect 415794 164898 415826 165134
rect 416062 164898 416146 165134
rect 416382 164898 416414 165134
rect 415794 129454 416414 164898
rect 415794 129218 415826 129454
rect 416062 129218 416146 129454
rect 416382 129218 416414 129454
rect 415794 129134 416414 129218
rect 415794 128898 415826 129134
rect 416062 128898 416146 129134
rect 416382 128898 416414 129134
rect 415794 93454 416414 128898
rect 415794 93218 415826 93454
rect 416062 93218 416146 93454
rect 416382 93218 416414 93454
rect 415794 93134 416414 93218
rect 415794 92898 415826 93134
rect 416062 92898 416146 93134
rect 416382 92898 416414 93134
rect 415794 57454 416414 92898
rect 415794 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 416414 57454
rect 415794 57134 416414 57218
rect 415794 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 416414 57134
rect 415794 21454 416414 56898
rect 415794 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 416414 21454
rect 415794 21134 416414 21218
rect 415794 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 416414 21134
rect 415794 -1306 416414 20898
rect 415794 -1542 415826 -1306
rect 416062 -1542 416146 -1306
rect 416382 -1542 416414 -1306
rect 415794 -1626 416414 -1542
rect 415794 -1862 415826 -1626
rect 416062 -1862 416146 -1626
rect 416382 -1862 416414 -1626
rect 415794 -1894 416414 -1862
rect 419514 169174 420134 198800
rect 419514 168938 419546 169174
rect 419782 168938 419866 169174
rect 420102 168938 420134 169174
rect 419514 168854 420134 168938
rect 419514 168618 419546 168854
rect 419782 168618 419866 168854
rect 420102 168618 420134 168854
rect 419514 133174 420134 168618
rect 419514 132938 419546 133174
rect 419782 132938 419866 133174
rect 420102 132938 420134 133174
rect 419514 132854 420134 132938
rect 419514 132618 419546 132854
rect 419782 132618 419866 132854
rect 420102 132618 420134 132854
rect 419514 97174 420134 132618
rect 419514 96938 419546 97174
rect 419782 96938 419866 97174
rect 420102 96938 420134 97174
rect 419514 96854 420134 96938
rect 419514 96618 419546 96854
rect 419782 96618 419866 96854
rect 420102 96618 420134 96854
rect 419514 61174 420134 96618
rect 419514 60938 419546 61174
rect 419782 60938 419866 61174
rect 420102 60938 420134 61174
rect 419514 60854 420134 60938
rect 419514 60618 419546 60854
rect 419782 60618 419866 60854
rect 420102 60618 420134 60854
rect 419514 25174 420134 60618
rect 419514 24938 419546 25174
rect 419782 24938 419866 25174
rect 420102 24938 420134 25174
rect 419514 24854 420134 24938
rect 419514 24618 419546 24854
rect 419782 24618 419866 24854
rect 420102 24618 420134 24854
rect 419514 -3226 420134 24618
rect 419514 -3462 419546 -3226
rect 419782 -3462 419866 -3226
rect 420102 -3462 420134 -3226
rect 419514 -3546 420134 -3462
rect 419514 -3782 419546 -3546
rect 419782 -3782 419866 -3546
rect 420102 -3782 420134 -3546
rect 419514 -3814 420134 -3782
rect 423234 172894 423854 208338
rect 423234 172658 423266 172894
rect 423502 172658 423586 172894
rect 423822 172658 423854 172894
rect 423234 172574 423854 172658
rect 423234 172338 423266 172574
rect 423502 172338 423586 172574
rect 423822 172338 423854 172574
rect 423234 136894 423854 172338
rect 423234 136658 423266 136894
rect 423502 136658 423586 136894
rect 423822 136658 423854 136894
rect 423234 136574 423854 136658
rect 423234 136338 423266 136574
rect 423502 136338 423586 136574
rect 423822 136338 423854 136574
rect 423234 100894 423854 136338
rect 423234 100658 423266 100894
rect 423502 100658 423586 100894
rect 423822 100658 423854 100894
rect 423234 100574 423854 100658
rect 423234 100338 423266 100574
rect 423502 100338 423586 100574
rect 423822 100338 423854 100574
rect 423234 64894 423854 100338
rect 423234 64658 423266 64894
rect 423502 64658 423586 64894
rect 423822 64658 423854 64894
rect 423234 64574 423854 64658
rect 423234 64338 423266 64574
rect 423502 64338 423586 64574
rect 423822 64338 423854 64574
rect 423234 28894 423854 64338
rect 423234 28658 423266 28894
rect 423502 28658 423586 28894
rect 423822 28658 423854 28894
rect 423234 28574 423854 28658
rect 423234 28338 423266 28574
rect 423502 28338 423586 28574
rect 423822 28338 423854 28574
rect 423234 -5146 423854 28338
rect 423234 -5382 423266 -5146
rect 423502 -5382 423586 -5146
rect 423822 -5382 423854 -5146
rect 423234 -5466 423854 -5382
rect 423234 -5702 423266 -5466
rect 423502 -5702 423586 -5466
rect 423822 -5702 423854 -5466
rect 423234 -5734 423854 -5702
rect 426954 680614 427574 711002
rect 444954 710598 445574 711590
rect 444954 710362 444986 710598
rect 445222 710362 445306 710598
rect 445542 710362 445574 710598
rect 444954 710278 445574 710362
rect 444954 710042 444986 710278
rect 445222 710042 445306 710278
rect 445542 710042 445574 710278
rect 441234 708678 441854 709670
rect 441234 708442 441266 708678
rect 441502 708442 441586 708678
rect 441822 708442 441854 708678
rect 441234 708358 441854 708442
rect 441234 708122 441266 708358
rect 441502 708122 441586 708358
rect 441822 708122 441854 708358
rect 437514 706758 438134 707750
rect 437514 706522 437546 706758
rect 437782 706522 437866 706758
rect 438102 706522 438134 706758
rect 437514 706438 438134 706522
rect 437514 706202 437546 706438
rect 437782 706202 437866 706438
rect 438102 706202 438134 706438
rect 426954 680378 426986 680614
rect 427222 680378 427306 680614
rect 427542 680378 427574 680614
rect 426954 680294 427574 680378
rect 426954 680058 426986 680294
rect 427222 680058 427306 680294
rect 427542 680058 427574 680294
rect 426954 644614 427574 680058
rect 426954 644378 426986 644614
rect 427222 644378 427306 644614
rect 427542 644378 427574 644614
rect 426954 644294 427574 644378
rect 426954 644058 426986 644294
rect 427222 644058 427306 644294
rect 427542 644058 427574 644294
rect 426954 608614 427574 644058
rect 426954 608378 426986 608614
rect 427222 608378 427306 608614
rect 427542 608378 427574 608614
rect 426954 608294 427574 608378
rect 426954 608058 426986 608294
rect 427222 608058 427306 608294
rect 427542 608058 427574 608294
rect 426954 572614 427574 608058
rect 426954 572378 426986 572614
rect 427222 572378 427306 572614
rect 427542 572378 427574 572614
rect 426954 572294 427574 572378
rect 426954 572058 426986 572294
rect 427222 572058 427306 572294
rect 427542 572058 427574 572294
rect 426954 536614 427574 572058
rect 426954 536378 426986 536614
rect 427222 536378 427306 536614
rect 427542 536378 427574 536614
rect 426954 536294 427574 536378
rect 426954 536058 426986 536294
rect 427222 536058 427306 536294
rect 427542 536058 427574 536294
rect 426954 500614 427574 536058
rect 426954 500378 426986 500614
rect 427222 500378 427306 500614
rect 427542 500378 427574 500614
rect 426954 500294 427574 500378
rect 426954 500058 426986 500294
rect 427222 500058 427306 500294
rect 427542 500058 427574 500294
rect 426954 464614 427574 500058
rect 426954 464378 426986 464614
rect 427222 464378 427306 464614
rect 427542 464378 427574 464614
rect 426954 464294 427574 464378
rect 426954 464058 426986 464294
rect 427222 464058 427306 464294
rect 427542 464058 427574 464294
rect 426954 428614 427574 464058
rect 426954 428378 426986 428614
rect 427222 428378 427306 428614
rect 427542 428378 427574 428614
rect 426954 428294 427574 428378
rect 426954 428058 426986 428294
rect 427222 428058 427306 428294
rect 427542 428058 427574 428294
rect 426954 392614 427574 428058
rect 426954 392378 426986 392614
rect 427222 392378 427306 392614
rect 427542 392378 427574 392614
rect 426954 392294 427574 392378
rect 426954 392058 426986 392294
rect 427222 392058 427306 392294
rect 427542 392058 427574 392294
rect 426954 356614 427574 392058
rect 426954 356378 426986 356614
rect 427222 356378 427306 356614
rect 427542 356378 427574 356614
rect 426954 356294 427574 356378
rect 426954 356058 426986 356294
rect 427222 356058 427306 356294
rect 427542 356058 427574 356294
rect 426954 320614 427574 356058
rect 426954 320378 426986 320614
rect 427222 320378 427306 320614
rect 427542 320378 427574 320614
rect 426954 320294 427574 320378
rect 426954 320058 426986 320294
rect 427222 320058 427306 320294
rect 427542 320058 427574 320294
rect 426954 284614 427574 320058
rect 426954 284378 426986 284614
rect 427222 284378 427306 284614
rect 427542 284378 427574 284614
rect 426954 284294 427574 284378
rect 426954 284058 426986 284294
rect 427222 284058 427306 284294
rect 427542 284058 427574 284294
rect 426954 248614 427574 284058
rect 426954 248378 426986 248614
rect 427222 248378 427306 248614
rect 427542 248378 427574 248614
rect 426954 248294 427574 248378
rect 426954 248058 426986 248294
rect 427222 248058 427306 248294
rect 427542 248058 427574 248294
rect 426954 212614 427574 248058
rect 426954 212378 426986 212614
rect 427222 212378 427306 212614
rect 427542 212378 427574 212614
rect 426954 212294 427574 212378
rect 426954 212058 426986 212294
rect 427222 212058 427306 212294
rect 427542 212058 427574 212294
rect 426954 176614 427574 212058
rect 426954 176378 426986 176614
rect 427222 176378 427306 176614
rect 427542 176378 427574 176614
rect 426954 176294 427574 176378
rect 426954 176058 426986 176294
rect 427222 176058 427306 176294
rect 427542 176058 427574 176294
rect 426954 140614 427574 176058
rect 426954 140378 426986 140614
rect 427222 140378 427306 140614
rect 427542 140378 427574 140614
rect 426954 140294 427574 140378
rect 426954 140058 426986 140294
rect 427222 140058 427306 140294
rect 427542 140058 427574 140294
rect 426954 104614 427574 140058
rect 426954 104378 426986 104614
rect 427222 104378 427306 104614
rect 427542 104378 427574 104614
rect 426954 104294 427574 104378
rect 426954 104058 426986 104294
rect 427222 104058 427306 104294
rect 427542 104058 427574 104294
rect 426954 68614 427574 104058
rect 426954 68378 426986 68614
rect 427222 68378 427306 68614
rect 427542 68378 427574 68614
rect 426954 68294 427574 68378
rect 426954 68058 426986 68294
rect 427222 68058 427306 68294
rect 427542 68058 427574 68294
rect 426954 32614 427574 68058
rect 426954 32378 426986 32614
rect 427222 32378 427306 32614
rect 427542 32378 427574 32614
rect 426954 32294 427574 32378
rect 426954 32058 426986 32294
rect 427222 32058 427306 32294
rect 427542 32058 427574 32294
rect 408954 -6342 408986 -6106
rect 409222 -6342 409306 -6106
rect 409542 -6342 409574 -6106
rect 408954 -6426 409574 -6342
rect 408954 -6662 408986 -6426
rect 409222 -6662 409306 -6426
rect 409542 -6662 409574 -6426
rect 408954 -7654 409574 -6662
rect 426954 -7066 427574 32058
rect 433794 704838 434414 705830
rect 433794 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 434414 704838
rect 433794 704518 434414 704602
rect 433794 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 434414 704518
rect 433794 687454 434414 704282
rect 433794 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 434414 687454
rect 433794 687134 434414 687218
rect 433794 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 434414 687134
rect 433794 651454 434414 686898
rect 433794 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 434414 651454
rect 433794 651134 434414 651218
rect 433794 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 434414 651134
rect 433794 615454 434414 650898
rect 433794 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 434414 615454
rect 433794 615134 434414 615218
rect 433794 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 434414 615134
rect 433794 579454 434414 614898
rect 433794 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 434414 579454
rect 433794 579134 434414 579218
rect 433794 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 434414 579134
rect 433794 543454 434414 578898
rect 433794 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 434414 543454
rect 433794 543134 434414 543218
rect 433794 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 434414 543134
rect 433794 507454 434414 542898
rect 433794 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 434414 507454
rect 433794 507134 434414 507218
rect 433794 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 434414 507134
rect 433794 471454 434414 506898
rect 433794 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 434414 471454
rect 433794 471134 434414 471218
rect 433794 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 434414 471134
rect 433794 435454 434414 470898
rect 433794 435218 433826 435454
rect 434062 435218 434146 435454
rect 434382 435218 434414 435454
rect 433794 435134 434414 435218
rect 433794 434898 433826 435134
rect 434062 434898 434146 435134
rect 434382 434898 434414 435134
rect 433794 399454 434414 434898
rect 433794 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 434414 399454
rect 433794 399134 434414 399218
rect 433794 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 434414 399134
rect 433794 363454 434414 398898
rect 433794 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 434414 363454
rect 433794 363134 434414 363218
rect 433794 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 434414 363134
rect 433794 327454 434414 362898
rect 433794 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 434414 327454
rect 433794 327134 434414 327218
rect 433794 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 434414 327134
rect 433794 291454 434414 326898
rect 433794 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 434414 291454
rect 433794 291134 434414 291218
rect 433794 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 434414 291134
rect 433794 255454 434414 290898
rect 433794 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 434414 255454
rect 433794 255134 434414 255218
rect 433794 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 434414 255134
rect 433794 219454 434414 254898
rect 433794 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 434414 219454
rect 433794 219134 434414 219218
rect 433794 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 434414 219134
rect 433794 183454 434414 218898
rect 433794 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 434414 183454
rect 433794 183134 434414 183218
rect 433794 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 434414 183134
rect 433794 147454 434414 182898
rect 433794 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 434414 147454
rect 433794 147134 434414 147218
rect 433794 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 434414 147134
rect 433794 111454 434414 146898
rect 433794 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 434414 111454
rect 433794 111134 434414 111218
rect 433794 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 434414 111134
rect 433794 75454 434414 110898
rect 433794 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 434414 75454
rect 433794 75134 434414 75218
rect 433794 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 434414 75134
rect 433794 39454 434414 74898
rect 433794 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 434414 39454
rect 433794 39134 434414 39218
rect 433794 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 434414 39134
rect 433794 3454 434414 38898
rect 433794 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 434414 3454
rect 433794 3134 434414 3218
rect 433794 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 434414 3134
rect 433794 -346 434414 2898
rect 433794 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 434414 -346
rect 433794 -666 434414 -582
rect 433794 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 434414 -666
rect 433794 -1894 434414 -902
rect 437514 691174 438134 706202
rect 437514 690938 437546 691174
rect 437782 690938 437866 691174
rect 438102 690938 438134 691174
rect 437514 690854 438134 690938
rect 437514 690618 437546 690854
rect 437782 690618 437866 690854
rect 438102 690618 438134 690854
rect 437514 655174 438134 690618
rect 437514 654938 437546 655174
rect 437782 654938 437866 655174
rect 438102 654938 438134 655174
rect 437514 654854 438134 654938
rect 437514 654618 437546 654854
rect 437782 654618 437866 654854
rect 438102 654618 438134 654854
rect 437514 619174 438134 654618
rect 437514 618938 437546 619174
rect 437782 618938 437866 619174
rect 438102 618938 438134 619174
rect 437514 618854 438134 618938
rect 437514 618618 437546 618854
rect 437782 618618 437866 618854
rect 438102 618618 438134 618854
rect 437514 583174 438134 618618
rect 437514 582938 437546 583174
rect 437782 582938 437866 583174
rect 438102 582938 438134 583174
rect 437514 582854 438134 582938
rect 437514 582618 437546 582854
rect 437782 582618 437866 582854
rect 438102 582618 438134 582854
rect 437514 547174 438134 582618
rect 437514 546938 437546 547174
rect 437782 546938 437866 547174
rect 438102 546938 438134 547174
rect 437514 546854 438134 546938
rect 437514 546618 437546 546854
rect 437782 546618 437866 546854
rect 438102 546618 438134 546854
rect 437514 511174 438134 546618
rect 437514 510938 437546 511174
rect 437782 510938 437866 511174
rect 438102 510938 438134 511174
rect 437514 510854 438134 510938
rect 437514 510618 437546 510854
rect 437782 510618 437866 510854
rect 438102 510618 438134 510854
rect 437514 475174 438134 510618
rect 437514 474938 437546 475174
rect 437782 474938 437866 475174
rect 438102 474938 438134 475174
rect 437514 474854 438134 474938
rect 437514 474618 437546 474854
rect 437782 474618 437866 474854
rect 438102 474618 438134 474854
rect 437514 439174 438134 474618
rect 437514 438938 437546 439174
rect 437782 438938 437866 439174
rect 438102 438938 438134 439174
rect 437514 438854 438134 438938
rect 437514 438618 437546 438854
rect 437782 438618 437866 438854
rect 438102 438618 438134 438854
rect 437514 403174 438134 438618
rect 437514 402938 437546 403174
rect 437782 402938 437866 403174
rect 438102 402938 438134 403174
rect 437514 402854 438134 402938
rect 437514 402618 437546 402854
rect 437782 402618 437866 402854
rect 438102 402618 438134 402854
rect 437514 367174 438134 402618
rect 437514 366938 437546 367174
rect 437782 366938 437866 367174
rect 438102 366938 438134 367174
rect 437514 366854 438134 366938
rect 437514 366618 437546 366854
rect 437782 366618 437866 366854
rect 438102 366618 438134 366854
rect 437514 331174 438134 366618
rect 437514 330938 437546 331174
rect 437782 330938 437866 331174
rect 438102 330938 438134 331174
rect 437514 330854 438134 330938
rect 437514 330618 437546 330854
rect 437782 330618 437866 330854
rect 438102 330618 438134 330854
rect 437514 295174 438134 330618
rect 437514 294938 437546 295174
rect 437782 294938 437866 295174
rect 438102 294938 438134 295174
rect 437514 294854 438134 294938
rect 437514 294618 437546 294854
rect 437782 294618 437866 294854
rect 438102 294618 438134 294854
rect 437514 259174 438134 294618
rect 437514 258938 437546 259174
rect 437782 258938 437866 259174
rect 438102 258938 438134 259174
rect 437514 258854 438134 258938
rect 437514 258618 437546 258854
rect 437782 258618 437866 258854
rect 438102 258618 438134 258854
rect 437514 223174 438134 258618
rect 437514 222938 437546 223174
rect 437782 222938 437866 223174
rect 438102 222938 438134 223174
rect 437514 222854 438134 222938
rect 437514 222618 437546 222854
rect 437782 222618 437866 222854
rect 438102 222618 438134 222854
rect 437514 187174 438134 222618
rect 437514 186938 437546 187174
rect 437782 186938 437866 187174
rect 438102 186938 438134 187174
rect 437514 186854 438134 186938
rect 437514 186618 437546 186854
rect 437782 186618 437866 186854
rect 438102 186618 438134 186854
rect 437514 151174 438134 186618
rect 437514 150938 437546 151174
rect 437782 150938 437866 151174
rect 438102 150938 438134 151174
rect 437514 150854 438134 150938
rect 437514 150618 437546 150854
rect 437782 150618 437866 150854
rect 438102 150618 438134 150854
rect 437514 115174 438134 150618
rect 437514 114938 437546 115174
rect 437782 114938 437866 115174
rect 438102 114938 438134 115174
rect 437514 114854 438134 114938
rect 437514 114618 437546 114854
rect 437782 114618 437866 114854
rect 438102 114618 438134 114854
rect 437514 79174 438134 114618
rect 437514 78938 437546 79174
rect 437782 78938 437866 79174
rect 438102 78938 438134 79174
rect 437514 78854 438134 78938
rect 437514 78618 437546 78854
rect 437782 78618 437866 78854
rect 438102 78618 438134 78854
rect 437514 43174 438134 78618
rect 437514 42938 437546 43174
rect 437782 42938 437866 43174
rect 438102 42938 438134 43174
rect 437514 42854 438134 42938
rect 437514 42618 437546 42854
rect 437782 42618 437866 42854
rect 438102 42618 438134 42854
rect 437514 7174 438134 42618
rect 437514 6938 437546 7174
rect 437782 6938 437866 7174
rect 438102 6938 438134 7174
rect 437514 6854 438134 6938
rect 437514 6618 437546 6854
rect 437782 6618 437866 6854
rect 438102 6618 438134 6854
rect 437514 -2266 438134 6618
rect 437514 -2502 437546 -2266
rect 437782 -2502 437866 -2266
rect 438102 -2502 438134 -2266
rect 437514 -2586 438134 -2502
rect 437514 -2822 437546 -2586
rect 437782 -2822 437866 -2586
rect 438102 -2822 438134 -2586
rect 437514 -3814 438134 -2822
rect 441234 694894 441854 708122
rect 441234 694658 441266 694894
rect 441502 694658 441586 694894
rect 441822 694658 441854 694894
rect 441234 694574 441854 694658
rect 441234 694338 441266 694574
rect 441502 694338 441586 694574
rect 441822 694338 441854 694574
rect 441234 658894 441854 694338
rect 441234 658658 441266 658894
rect 441502 658658 441586 658894
rect 441822 658658 441854 658894
rect 441234 658574 441854 658658
rect 441234 658338 441266 658574
rect 441502 658338 441586 658574
rect 441822 658338 441854 658574
rect 441234 622894 441854 658338
rect 441234 622658 441266 622894
rect 441502 622658 441586 622894
rect 441822 622658 441854 622894
rect 441234 622574 441854 622658
rect 441234 622338 441266 622574
rect 441502 622338 441586 622574
rect 441822 622338 441854 622574
rect 441234 586894 441854 622338
rect 441234 586658 441266 586894
rect 441502 586658 441586 586894
rect 441822 586658 441854 586894
rect 441234 586574 441854 586658
rect 441234 586338 441266 586574
rect 441502 586338 441586 586574
rect 441822 586338 441854 586574
rect 441234 550894 441854 586338
rect 441234 550658 441266 550894
rect 441502 550658 441586 550894
rect 441822 550658 441854 550894
rect 441234 550574 441854 550658
rect 441234 550338 441266 550574
rect 441502 550338 441586 550574
rect 441822 550338 441854 550574
rect 441234 514894 441854 550338
rect 441234 514658 441266 514894
rect 441502 514658 441586 514894
rect 441822 514658 441854 514894
rect 441234 514574 441854 514658
rect 441234 514338 441266 514574
rect 441502 514338 441586 514574
rect 441822 514338 441854 514574
rect 441234 478894 441854 514338
rect 441234 478658 441266 478894
rect 441502 478658 441586 478894
rect 441822 478658 441854 478894
rect 441234 478574 441854 478658
rect 441234 478338 441266 478574
rect 441502 478338 441586 478574
rect 441822 478338 441854 478574
rect 441234 442894 441854 478338
rect 441234 442658 441266 442894
rect 441502 442658 441586 442894
rect 441822 442658 441854 442894
rect 441234 442574 441854 442658
rect 441234 442338 441266 442574
rect 441502 442338 441586 442574
rect 441822 442338 441854 442574
rect 441234 406894 441854 442338
rect 441234 406658 441266 406894
rect 441502 406658 441586 406894
rect 441822 406658 441854 406894
rect 441234 406574 441854 406658
rect 441234 406338 441266 406574
rect 441502 406338 441586 406574
rect 441822 406338 441854 406574
rect 441234 370894 441854 406338
rect 441234 370658 441266 370894
rect 441502 370658 441586 370894
rect 441822 370658 441854 370894
rect 441234 370574 441854 370658
rect 441234 370338 441266 370574
rect 441502 370338 441586 370574
rect 441822 370338 441854 370574
rect 441234 334894 441854 370338
rect 441234 334658 441266 334894
rect 441502 334658 441586 334894
rect 441822 334658 441854 334894
rect 441234 334574 441854 334658
rect 441234 334338 441266 334574
rect 441502 334338 441586 334574
rect 441822 334338 441854 334574
rect 441234 298894 441854 334338
rect 441234 298658 441266 298894
rect 441502 298658 441586 298894
rect 441822 298658 441854 298894
rect 441234 298574 441854 298658
rect 441234 298338 441266 298574
rect 441502 298338 441586 298574
rect 441822 298338 441854 298574
rect 441234 262894 441854 298338
rect 441234 262658 441266 262894
rect 441502 262658 441586 262894
rect 441822 262658 441854 262894
rect 441234 262574 441854 262658
rect 441234 262338 441266 262574
rect 441502 262338 441586 262574
rect 441822 262338 441854 262574
rect 441234 226894 441854 262338
rect 441234 226658 441266 226894
rect 441502 226658 441586 226894
rect 441822 226658 441854 226894
rect 441234 226574 441854 226658
rect 441234 226338 441266 226574
rect 441502 226338 441586 226574
rect 441822 226338 441854 226574
rect 441234 190894 441854 226338
rect 441234 190658 441266 190894
rect 441502 190658 441586 190894
rect 441822 190658 441854 190894
rect 441234 190574 441854 190658
rect 441234 190338 441266 190574
rect 441502 190338 441586 190574
rect 441822 190338 441854 190574
rect 441234 154894 441854 190338
rect 441234 154658 441266 154894
rect 441502 154658 441586 154894
rect 441822 154658 441854 154894
rect 441234 154574 441854 154658
rect 441234 154338 441266 154574
rect 441502 154338 441586 154574
rect 441822 154338 441854 154574
rect 441234 118894 441854 154338
rect 441234 118658 441266 118894
rect 441502 118658 441586 118894
rect 441822 118658 441854 118894
rect 441234 118574 441854 118658
rect 441234 118338 441266 118574
rect 441502 118338 441586 118574
rect 441822 118338 441854 118574
rect 441234 82894 441854 118338
rect 441234 82658 441266 82894
rect 441502 82658 441586 82894
rect 441822 82658 441854 82894
rect 441234 82574 441854 82658
rect 441234 82338 441266 82574
rect 441502 82338 441586 82574
rect 441822 82338 441854 82574
rect 441234 46894 441854 82338
rect 441234 46658 441266 46894
rect 441502 46658 441586 46894
rect 441822 46658 441854 46894
rect 441234 46574 441854 46658
rect 441234 46338 441266 46574
rect 441502 46338 441586 46574
rect 441822 46338 441854 46574
rect 441234 10894 441854 46338
rect 441234 10658 441266 10894
rect 441502 10658 441586 10894
rect 441822 10658 441854 10894
rect 441234 10574 441854 10658
rect 441234 10338 441266 10574
rect 441502 10338 441586 10574
rect 441822 10338 441854 10574
rect 441234 -4186 441854 10338
rect 441234 -4422 441266 -4186
rect 441502 -4422 441586 -4186
rect 441822 -4422 441854 -4186
rect 441234 -4506 441854 -4422
rect 441234 -4742 441266 -4506
rect 441502 -4742 441586 -4506
rect 441822 -4742 441854 -4506
rect 441234 -5734 441854 -4742
rect 444954 698614 445574 710042
rect 462954 711558 463574 711590
rect 462954 711322 462986 711558
rect 463222 711322 463306 711558
rect 463542 711322 463574 711558
rect 462954 711238 463574 711322
rect 462954 711002 462986 711238
rect 463222 711002 463306 711238
rect 463542 711002 463574 711238
rect 459234 709638 459854 709670
rect 459234 709402 459266 709638
rect 459502 709402 459586 709638
rect 459822 709402 459854 709638
rect 459234 709318 459854 709402
rect 459234 709082 459266 709318
rect 459502 709082 459586 709318
rect 459822 709082 459854 709318
rect 455514 707718 456134 707750
rect 455514 707482 455546 707718
rect 455782 707482 455866 707718
rect 456102 707482 456134 707718
rect 455514 707398 456134 707482
rect 455514 707162 455546 707398
rect 455782 707162 455866 707398
rect 456102 707162 456134 707398
rect 444954 698378 444986 698614
rect 445222 698378 445306 698614
rect 445542 698378 445574 698614
rect 444954 698294 445574 698378
rect 444954 698058 444986 698294
rect 445222 698058 445306 698294
rect 445542 698058 445574 698294
rect 444954 662614 445574 698058
rect 444954 662378 444986 662614
rect 445222 662378 445306 662614
rect 445542 662378 445574 662614
rect 444954 662294 445574 662378
rect 444954 662058 444986 662294
rect 445222 662058 445306 662294
rect 445542 662058 445574 662294
rect 444954 626614 445574 662058
rect 444954 626378 444986 626614
rect 445222 626378 445306 626614
rect 445542 626378 445574 626614
rect 444954 626294 445574 626378
rect 444954 626058 444986 626294
rect 445222 626058 445306 626294
rect 445542 626058 445574 626294
rect 444954 590614 445574 626058
rect 444954 590378 444986 590614
rect 445222 590378 445306 590614
rect 445542 590378 445574 590614
rect 444954 590294 445574 590378
rect 444954 590058 444986 590294
rect 445222 590058 445306 590294
rect 445542 590058 445574 590294
rect 444954 554614 445574 590058
rect 444954 554378 444986 554614
rect 445222 554378 445306 554614
rect 445542 554378 445574 554614
rect 444954 554294 445574 554378
rect 444954 554058 444986 554294
rect 445222 554058 445306 554294
rect 445542 554058 445574 554294
rect 444954 518614 445574 554058
rect 444954 518378 444986 518614
rect 445222 518378 445306 518614
rect 445542 518378 445574 518614
rect 444954 518294 445574 518378
rect 444954 518058 444986 518294
rect 445222 518058 445306 518294
rect 445542 518058 445574 518294
rect 444954 482614 445574 518058
rect 444954 482378 444986 482614
rect 445222 482378 445306 482614
rect 445542 482378 445574 482614
rect 444954 482294 445574 482378
rect 444954 482058 444986 482294
rect 445222 482058 445306 482294
rect 445542 482058 445574 482294
rect 444954 446614 445574 482058
rect 444954 446378 444986 446614
rect 445222 446378 445306 446614
rect 445542 446378 445574 446614
rect 444954 446294 445574 446378
rect 444954 446058 444986 446294
rect 445222 446058 445306 446294
rect 445542 446058 445574 446294
rect 444954 410614 445574 446058
rect 444954 410378 444986 410614
rect 445222 410378 445306 410614
rect 445542 410378 445574 410614
rect 444954 410294 445574 410378
rect 444954 410058 444986 410294
rect 445222 410058 445306 410294
rect 445542 410058 445574 410294
rect 444954 374614 445574 410058
rect 444954 374378 444986 374614
rect 445222 374378 445306 374614
rect 445542 374378 445574 374614
rect 444954 374294 445574 374378
rect 444954 374058 444986 374294
rect 445222 374058 445306 374294
rect 445542 374058 445574 374294
rect 444954 338614 445574 374058
rect 444954 338378 444986 338614
rect 445222 338378 445306 338614
rect 445542 338378 445574 338614
rect 444954 338294 445574 338378
rect 444954 338058 444986 338294
rect 445222 338058 445306 338294
rect 445542 338058 445574 338294
rect 444954 302614 445574 338058
rect 444954 302378 444986 302614
rect 445222 302378 445306 302614
rect 445542 302378 445574 302614
rect 444954 302294 445574 302378
rect 444954 302058 444986 302294
rect 445222 302058 445306 302294
rect 445542 302058 445574 302294
rect 444954 266614 445574 302058
rect 444954 266378 444986 266614
rect 445222 266378 445306 266614
rect 445542 266378 445574 266614
rect 444954 266294 445574 266378
rect 444954 266058 444986 266294
rect 445222 266058 445306 266294
rect 445542 266058 445574 266294
rect 444954 230614 445574 266058
rect 444954 230378 444986 230614
rect 445222 230378 445306 230614
rect 445542 230378 445574 230614
rect 444954 230294 445574 230378
rect 444954 230058 444986 230294
rect 445222 230058 445306 230294
rect 445542 230058 445574 230294
rect 444954 194614 445574 230058
rect 444954 194378 444986 194614
rect 445222 194378 445306 194614
rect 445542 194378 445574 194614
rect 444954 194294 445574 194378
rect 444954 194058 444986 194294
rect 445222 194058 445306 194294
rect 445542 194058 445574 194294
rect 444954 158614 445574 194058
rect 444954 158378 444986 158614
rect 445222 158378 445306 158614
rect 445542 158378 445574 158614
rect 444954 158294 445574 158378
rect 444954 158058 444986 158294
rect 445222 158058 445306 158294
rect 445542 158058 445574 158294
rect 444954 122614 445574 158058
rect 444954 122378 444986 122614
rect 445222 122378 445306 122614
rect 445542 122378 445574 122614
rect 444954 122294 445574 122378
rect 444954 122058 444986 122294
rect 445222 122058 445306 122294
rect 445542 122058 445574 122294
rect 444954 86614 445574 122058
rect 444954 86378 444986 86614
rect 445222 86378 445306 86614
rect 445542 86378 445574 86614
rect 444954 86294 445574 86378
rect 444954 86058 444986 86294
rect 445222 86058 445306 86294
rect 445542 86058 445574 86294
rect 444954 50614 445574 86058
rect 444954 50378 444986 50614
rect 445222 50378 445306 50614
rect 445542 50378 445574 50614
rect 444954 50294 445574 50378
rect 444954 50058 444986 50294
rect 445222 50058 445306 50294
rect 445542 50058 445574 50294
rect 444954 14614 445574 50058
rect 444954 14378 444986 14614
rect 445222 14378 445306 14614
rect 445542 14378 445574 14614
rect 444954 14294 445574 14378
rect 444954 14058 444986 14294
rect 445222 14058 445306 14294
rect 445542 14058 445574 14294
rect 426954 -7302 426986 -7066
rect 427222 -7302 427306 -7066
rect 427542 -7302 427574 -7066
rect 426954 -7386 427574 -7302
rect 426954 -7622 426986 -7386
rect 427222 -7622 427306 -7386
rect 427542 -7622 427574 -7386
rect 426954 -7654 427574 -7622
rect 444954 -6106 445574 14058
rect 451794 705798 452414 705830
rect 451794 705562 451826 705798
rect 452062 705562 452146 705798
rect 452382 705562 452414 705798
rect 451794 705478 452414 705562
rect 451794 705242 451826 705478
rect 452062 705242 452146 705478
rect 452382 705242 452414 705478
rect 451794 669454 452414 705242
rect 451794 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 452414 669454
rect 451794 669134 452414 669218
rect 451794 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 452414 669134
rect 451794 633454 452414 668898
rect 451794 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 452414 633454
rect 451794 633134 452414 633218
rect 451794 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 452414 633134
rect 451794 597454 452414 632898
rect 451794 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 452414 597454
rect 451794 597134 452414 597218
rect 451794 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 452414 597134
rect 451794 561454 452414 596898
rect 451794 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 452414 561454
rect 451794 561134 452414 561218
rect 451794 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 452414 561134
rect 451794 525454 452414 560898
rect 451794 525218 451826 525454
rect 452062 525218 452146 525454
rect 452382 525218 452414 525454
rect 451794 525134 452414 525218
rect 451794 524898 451826 525134
rect 452062 524898 452146 525134
rect 452382 524898 452414 525134
rect 451794 489454 452414 524898
rect 451794 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 452414 489454
rect 451794 489134 452414 489218
rect 451794 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 452414 489134
rect 451794 453454 452414 488898
rect 451794 453218 451826 453454
rect 452062 453218 452146 453454
rect 452382 453218 452414 453454
rect 451794 453134 452414 453218
rect 451794 452898 451826 453134
rect 452062 452898 452146 453134
rect 452382 452898 452414 453134
rect 451794 417454 452414 452898
rect 451794 417218 451826 417454
rect 452062 417218 452146 417454
rect 452382 417218 452414 417454
rect 451794 417134 452414 417218
rect 451794 416898 451826 417134
rect 452062 416898 452146 417134
rect 452382 416898 452414 417134
rect 451794 381454 452414 416898
rect 451794 381218 451826 381454
rect 452062 381218 452146 381454
rect 452382 381218 452414 381454
rect 451794 381134 452414 381218
rect 451794 380898 451826 381134
rect 452062 380898 452146 381134
rect 452382 380898 452414 381134
rect 451794 345454 452414 380898
rect 451794 345218 451826 345454
rect 452062 345218 452146 345454
rect 452382 345218 452414 345454
rect 451794 345134 452414 345218
rect 451794 344898 451826 345134
rect 452062 344898 452146 345134
rect 452382 344898 452414 345134
rect 451794 309454 452414 344898
rect 451794 309218 451826 309454
rect 452062 309218 452146 309454
rect 452382 309218 452414 309454
rect 451794 309134 452414 309218
rect 451794 308898 451826 309134
rect 452062 308898 452146 309134
rect 452382 308898 452414 309134
rect 451794 273454 452414 308898
rect 451794 273218 451826 273454
rect 452062 273218 452146 273454
rect 452382 273218 452414 273454
rect 451794 273134 452414 273218
rect 451794 272898 451826 273134
rect 452062 272898 452146 273134
rect 452382 272898 452414 273134
rect 451794 237454 452414 272898
rect 451794 237218 451826 237454
rect 452062 237218 452146 237454
rect 452382 237218 452414 237454
rect 451794 237134 452414 237218
rect 451794 236898 451826 237134
rect 452062 236898 452146 237134
rect 452382 236898 452414 237134
rect 451794 201454 452414 236898
rect 451794 201218 451826 201454
rect 452062 201218 452146 201454
rect 452382 201218 452414 201454
rect 451794 201134 452414 201218
rect 451794 200898 451826 201134
rect 452062 200898 452146 201134
rect 452382 200898 452414 201134
rect 451794 165454 452414 200898
rect 451794 165218 451826 165454
rect 452062 165218 452146 165454
rect 452382 165218 452414 165454
rect 451794 165134 452414 165218
rect 451794 164898 451826 165134
rect 452062 164898 452146 165134
rect 452382 164898 452414 165134
rect 451794 129454 452414 164898
rect 451794 129218 451826 129454
rect 452062 129218 452146 129454
rect 452382 129218 452414 129454
rect 451794 129134 452414 129218
rect 451794 128898 451826 129134
rect 452062 128898 452146 129134
rect 452382 128898 452414 129134
rect 451794 93454 452414 128898
rect 451794 93218 451826 93454
rect 452062 93218 452146 93454
rect 452382 93218 452414 93454
rect 451794 93134 452414 93218
rect 451794 92898 451826 93134
rect 452062 92898 452146 93134
rect 452382 92898 452414 93134
rect 451794 57454 452414 92898
rect 451794 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 452414 57454
rect 451794 57134 452414 57218
rect 451794 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 452414 57134
rect 451794 21454 452414 56898
rect 451794 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 452414 21454
rect 451794 21134 452414 21218
rect 451794 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 452414 21134
rect 451794 -1306 452414 20898
rect 451794 -1542 451826 -1306
rect 452062 -1542 452146 -1306
rect 452382 -1542 452414 -1306
rect 451794 -1626 452414 -1542
rect 451794 -1862 451826 -1626
rect 452062 -1862 452146 -1626
rect 452382 -1862 452414 -1626
rect 451794 -1894 452414 -1862
rect 455514 673174 456134 707162
rect 455514 672938 455546 673174
rect 455782 672938 455866 673174
rect 456102 672938 456134 673174
rect 455514 672854 456134 672938
rect 455514 672618 455546 672854
rect 455782 672618 455866 672854
rect 456102 672618 456134 672854
rect 455514 637174 456134 672618
rect 455514 636938 455546 637174
rect 455782 636938 455866 637174
rect 456102 636938 456134 637174
rect 455514 636854 456134 636938
rect 455514 636618 455546 636854
rect 455782 636618 455866 636854
rect 456102 636618 456134 636854
rect 455514 601174 456134 636618
rect 455514 600938 455546 601174
rect 455782 600938 455866 601174
rect 456102 600938 456134 601174
rect 455514 600854 456134 600938
rect 455514 600618 455546 600854
rect 455782 600618 455866 600854
rect 456102 600618 456134 600854
rect 455514 565174 456134 600618
rect 455514 564938 455546 565174
rect 455782 564938 455866 565174
rect 456102 564938 456134 565174
rect 455514 564854 456134 564938
rect 455514 564618 455546 564854
rect 455782 564618 455866 564854
rect 456102 564618 456134 564854
rect 455514 529174 456134 564618
rect 455514 528938 455546 529174
rect 455782 528938 455866 529174
rect 456102 528938 456134 529174
rect 455514 528854 456134 528938
rect 455514 528618 455546 528854
rect 455782 528618 455866 528854
rect 456102 528618 456134 528854
rect 455514 493174 456134 528618
rect 455514 492938 455546 493174
rect 455782 492938 455866 493174
rect 456102 492938 456134 493174
rect 455514 492854 456134 492938
rect 455514 492618 455546 492854
rect 455782 492618 455866 492854
rect 456102 492618 456134 492854
rect 455514 457174 456134 492618
rect 455514 456938 455546 457174
rect 455782 456938 455866 457174
rect 456102 456938 456134 457174
rect 455514 456854 456134 456938
rect 455514 456618 455546 456854
rect 455782 456618 455866 456854
rect 456102 456618 456134 456854
rect 455514 421174 456134 456618
rect 455514 420938 455546 421174
rect 455782 420938 455866 421174
rect 456102 420938 456134 421174
rect 455514 420854 456134 420938
rect 455514 420618 455546 420854
rect 455782 420618 455866 420854
rect 456102 420618 456134 420854
rect 455514 385174 456134 420618
rect 455514 384938 455546 385174
rect 455782 384938 455866 385174
rect 456102 384938 456134 385174
rect 455514 384854 456134 384938
rect 455514 384618 455546 384854
rect 455782 384618 455866 384854
rect 456102 384618 456134 384854
rect 455514 349174 456134 384618
rect 455514 348938 455546 349174
rect 455782 348938 455866 349174
rect 456102 348938 456134 349174
rect 455514 348854 456134 348938
rect 455514 348618 455546 348854
rect 455782 348618 455866 348854
rect 456102 348618 456134 348854
rect 455514 313174 456134 348618
rect 455514 312938 455546 313174
rect 455782 312938 455866 313174
rect 456102 312938 456134 313174
rect 455514 312854 456134 312938
rect 455514 312618 455546 312854
rect 455782 312618 455866 312854
rect 456102 312618 456134 312854
rect 455514 277174 456134 312618
rect 455514 276938 455546 277174
rect 455782 276938 455866 277174
rect 456102 276938 456134 277174
rect 455514 276854 456134 276938
rect 455514 276618 455546 276854
rect 455782 276618 455866 276854
rect 456102 276618 456134 276854
rect 455514 241174 456134 276618
rect 455514 240938 455546 241174
rect 455782 240938 455866 241174
rect 456102 240938 456134 241174
rect 455514 240854 456134 240938
rect 455514 240618 455546 240854
rect 455782 240618 455866 240854
rect 456102 240618 456134 240854
rect 455514 205174 456134 240618
rect 455514 204938 455546 205174
rect 455782 204938 455866 205174
rect 456102 204938 456134 205174
rect 455514 204854 456134 204938
rect 455514 204618 455546 204854
rect 455782 204618 455866 204854
rect 456102 204618 456134 204854
rect 455514 169174 456134 204618
rect 455514 168938 455546 169174
rect 455782 168938 455866 169174
rect 456102 168938 456134 169174
rect 455514 168854 456134 168938
rect 455514 168618 455546 168854
rect 455782 168618 455866 168854
rect 456102 168618 456134 168854
rect 455514 133174 456134 168618
rect 455514 132938 455546 133174
rect 455782 132938 455866 133174
rect 456102 132938 456134 133174
rect 455514 132854 456134 132938
rect 455514 132618 455546 132854
rect 455782 132618 455866 132854
rect 456102 132618 456134 132854
rect 455514 97174 456134 132618
rect 455514 96938 455546 97174
rect 455782 96938 455866 97174
rect 456102 96938 456134 97174
rect 455514 96854 456134 96938
rect 455514 96618 455546 96854
rect 455782 96618 455866 96854
rect 456102 96618 456134 96854
rect 455514 61174 456134 96618
rect 455514 60938 455546 61174
rect 455782 60938 455866 61174
rect 456102 60938 456134 61174
rect 455514 60854 456134 60938
rect 455514 60618 455546 60854
rect 455782 60618 455866 60854
rect 456102 60618 456134 60854
rect 455514 25174 456134 60618
rect 455514 24938 455546 25174
rect 455782 24938 455866 25174
rect 456102 24938 456134 25174
rect 455514 24854 456134 24938
rect 455514 24618 455546 24854
rect 455782 24618 455866 24854
rect 456102 24618 456134 24854
rect 455514 -3226 456134 24618
rect 455514 -3462 455546 -3226
rect 455782 -3462 455866 -3226
rect 456102 -3462 456134 -3226
rect 455514 -3546 456134 -3462
rect 455514 -3782 455546 -3546
rect 455782 -3782 455866 -3546
rect 456102 -3782 456134 -3546
rect 455514 -3814 456134 -3782
rect 459234 676894 459854 709082
rect 459234 676658 459266 676894
rect 459502 676658 459586 676894
rect 459822 676658 459854 676894
rect 459234 676574 459854 676658
rect 459234 676338 459266 676574
rect 459502 676338 459586 676574
rect 459822 676338 459854 676574
rect 459234 640894 459854 676338
rect 459234 640658 459266 640894
rect 459502 640658 459586 640894
rect 459822 640658 459854 640894
rect 459234 640574 459854 640658
rect 459234 640338 459266 640574
rect 459502 640338 459586 640574
rect 459822 640338 459854 640574
rect 459234 604894 459854 640338
rect 459234 604658 459266 604894
rect 459502 604658 459586 604894
rect 459822 604658 459854 604894
rect 459234 604574 459854 604658
rect 459234 604338 459266 604574
rect 459502 604338 459586 604574
rect 459822 604338 459854 604574
rect 459234 568894 459854 604338
rect 459234 568658 459266 568894
rect 459502 568658 459586 568894
rect 459822 568658 459854 568894
rect 459234 568574 459854 568658
rect 459234 568338 459266 568574
rect 459502 568338 459586 568574
rect 459822 568338 459854 568574
rect 459234 532894 459854 568338
rect 459234 532658 459266 532894
rect 459502 532658 459586 532894
rect 459822 532658 459854 532894
rect 459234 532574 459854 532658
rect 459234 532338 459266 532574
rect 459502 532338 459586 532574
rect 459822 532338 459854 532574
rect 459234 496894 459854 532338
rect 459234 496658 459266 496894
rect 459502 496658 459586 496894
rect 459822 496658 459854 496894
rect 459234 496574 459854 496658
rect 459234 496338 459266 496574
rect 459502 496338 459586 496574
rect 459822 496338 459854 496574
rect 459234 460894 459854 496338
rect 459234 460658 459266 460894
rect 459502 460658 459586 460894
rect 459822 460658 459854 460894
rect 459234 460574 459854 460658
rect 459234 460338 459266 460574
rect 459502 460338 459586 460574
rect 459822 460338 459854 460574
rect 459234 424894 459854 460338
rect 459234 424658 459266 424894
rect 459502 424658 459586 424894
rect 459822 424658 459854 424894
rect 459234 424574 459854 424658
rect 459234 424338 459266 424574
rect 459502 424338 459586 424574
rect 459822 424338 459854 424574
rect 459234 388894 459854 424338
rect 459234 388658 459266 388894
rect 459502 388658 459586 388894
rect 459822 388658 459854 388894
rect 459234 388574 459854 388658
rect 459234 388338 459266 388574
rect 459502 388338 459586 388574
rect 459822 388338 459854 388574
rect 459234 352894 459854 388338
rect 459234 352658 459266 352894
rect 459502 352658 459586 352894
rect 459822 352658 459854 352894
rect 459234 352574 459854 352658
rect 459234 352338 459266 352574
rect 459502 352338 459586 352574
rect 459822 352338 459854 352574
rect 459234 316894 459854 352338
rect 459234 316658 459266 316894
rect 459502 316658 459586 316894
rect 459822 316658 459854 316894
rect 459234 316574 459854 316658
rect 459234 316338 459266 316574
rect 459502 316338 459586 316574
rect 459822 316338 459854 316574
rect 459234 280894 459854 316338
rect 459234 280658 459266 280894
rect 459502 280658 459586 280894
rect 459822 280658 459854 280894
rect 459234 280574 459854 280658
rect 459234 280338 459266 280574
rect 459502 280338 459586 280574
rect 459822 280338 459854 280574
rect 459234 244894 459854 280338
rect 459234 244658 459266 244894
rect 459502 244658 459586 244894
rect 459822 244658 459854 244894
rect 459234 244574 459854 244658
rect 459234 244338 459266 244574
rect 459502 244338 459586 244574
rect 459822 244338 459854 244574
rect 459234 208894 459854 244338
rect 459234 208658 459266 208894
rect 459502 208658 459586 208894
rect 459822 208658 459854 208894
rect 459234 208574 459854 208658
rect 459234 208338 459266 208574
rect 459502 208338 459586 208574
rect 459822 208338 459854 208574
rect 459234 172894 459854 208338
rect 459234 172658 459266 172894
rect 459502 172658 459586 172894
rect 459822 172658 459854 172894
rect 459234 172574 459854 172658
rect 459234 172338 459266 172574
rect 459502 172338 459586 172574
rect 459822 172338 459854 172574
rect 459234 136894 459854 172338
rect 459234 136658 459266 136894
rect 459502 136658 459586 136894
rect 459822 136658 459854 136894
rect 459234 136574 459854 136658
rect 459234 136338 459266 136574
rect 459502 136338 459586 136574
rect 459822 136338 459854 136574
rect 459234 100894 459854 136338
rect 459234 100658 459266 100894
rect 459502 100658 459586 100894
rect 459822 100658 459854 100894
rect 459234 100574 459854 100658
rect 459234 100338 459266 100574
rect 459502 100338 459586 100574
rect 459822 100338 459854 100574
rect 459234 64894 459854 100338
rect 459234 64658 459266 64894
rect 459502 64658 459586 64894
rect 459822 64658 459854 64894
rect 459234 64574 459854 64658
rect 459234 64338 459266 64574
rect 459502 64338 459586 64574
rect 459822 64338 459854 64574
rect 459234 28894 459854 64338
rect 459234 28658 459266 28894
rect 459502 28658 459586 28894
rect 459822 28658 459854 28894
rect 459234 28574 459854 28658
rect 459234 28338 459266 28574
rect 459502 28338 459586 28574
rect 459822 28338 459854 28574
rect 459234 -5146 459854 28338
rect 459234 -5382 459266 -5146
rect 459502 -5382 459586 -5146
rect 459822 -5382 459854 -5146
rect 459234 -5466 459854 -5382
rect 459234 -5702 459266 -5466
rect 459502 -5702 459586 -5466
rect 459822 -5702 459854 -5466
rect 459234 -5734 459854 -5702
rect 462954 680614 463574 711002
rect 480954 710598 481574 711590
rect 480954 710362 480986 710598
rect 481222 710362 481306 710598
rect 481542 710362 481574 710598
rect 480954 710278 481574 710362
rect 480954 710042 480986 710278
rect 481222 710042 481306 710278
rect 481542 710042 481574 710278
rect 477234 708678 477854 709670
rect 477234 708442 477266 708678
rect 477502 708442 477586 708678
rect 477822 708442 477854 708678
rect 477234 708358 477854 708442
rect 477234 708122 477266 708358
rect 477502 708122 477586 708358
rect 477822 708122 477854 708358
rect 473514 706758 474134 707750
rect 473514 706522 473546 706758
rect 473782 706522 473866 706758
rect 474102 706522 474134 706758
rect 473514 706438 474134 706522
rect 473514 706202 473546 706438
rect 473782 706202 473866 706438
rect 474102 706202 474134 706438
rect 462954 680378 462986 680614
rect 463222 680378 463306 680614
rect 463542 680378 463574 680614
rect 462954 680294 463574 680378
rect 462954 680058 462986 680294
rect 463222 680058 463306 680294
rect 463542 680058 463574 680294
rect 462954 644614 463574 680058
rect 462954 644378 462986 644614
rect 463222 644378 463306 644614
rect 463542 644378 463574 644614
rect 462954 644294 463574 644378
rect 462954 644058 462986 644294
rect 463222 644058 463306 644294
rect 463542 644058 463574 644294
rect 462954 608614 463574 644058
rect 462954 608378 462986 608614
rect 463222 608378 463306 608614
rect 463542 608378 463574 608614
rect 462954 608294 463574 608378
rect 462954 608058 462986 608294
rect 463222 608058 463306 608294
rect 463542 608058 463574 608294
rect 462954 572614 463574 608058
rect 462954 572378 462986 572614
rect 463222 572378 463306 572614
rect 463542 572378 463574 572614
rect 462954 572294 463574 572378
rect 462954 572058 462986 572294
rect 463222 572058 463306 572294
rect 463542 572058 463574 572294
rect 462954 536614 463574 572058
rect 462954 536378 462986 536614
rect 463222 536378 463306 536614
rect 463542 536378 463574 536614
rect 462954 536294 463574 536378
rect 462954 536058 462986 536294
rect 463222 536058 463306 536294
rect 463542 536058 463574 536294
rect 462954 500614 463574 536058
rect 462954 500378 462986 500614
rect 463222 500378 463306 500614
rect 463542 500378 463574 500614
rect 462954 500294 463574 500378
rect 462954 500058 462986 500294
rect 463222 500058 463306 500294
rect 463542 500058 463574 500294
rect 462954 464614 463574 500058
rect 462954 464378 462986 464614
rect 463222 464378 463306 464614
rect 463542 464378 463574 464614
rect 462954 464294 463574 464378
rect 462954 464058 462986 464294
rect 463222 464058 463306 464294
rect 463542 464058 463574 464294
rect 462954 428614 463574 464058
rect 462954 428378 462986 428614
rect 463222 428378 463306 428614
rect 463542 428378 463574 428614
rect 462954 428294 463574 428378
rect 462954 428058 462986 428294
rect 463222 428058 463306 428294
rect 463542 428058 463574 428294
rect 462954 392614 463574 428058
rect 462954 392378 462986 392614
rect 463222 392378 463306 392614
rect 463542 392378 463574 392614
rect 462954 392294 463574 392378
rect 462954 392058 462986 392294
rect 463222 392058 463306 392294
rect 463542 392058 463574 392294
rect 462954 356614 463574 392058
rect 462954 356378 462986 356614
rect 463222 356378 463306 356614
rect 463542 356378 463574 356614
rect 462954 356294 463574 356378
rect 462954 356058 462986 356294
rect 463222 356058 463306 356294
rect 463542 356058 463574 356294
rect 462954 320614 463574 356058
rect 462954 320378 462986 320614
rect 463222 320378 463306 320614
rect 463542 320378 463574 320614
rect 462954 320294 463574 320378
rect 462954 320058 462986 320294
rect 463222 320058 463306 320294
rect 463542 320058 463574 320294
rect 462954 284614 463574 320058
rect 462954 284378 462986 284614
rect 463222 284378 463306 284614
rect 463542 284378 463574 284614
rect 462954 284294 463574 284378
rect 462954 284058 462986 284294
rect 463222 284058 463306 284294
rect 463542 284058 463574 284294
rect 462954 248614 463574 284058
rect 462954 248378 462986 248614
rect 463222 248378 463306 248614
rect 463542 248378 463574 248614
rect 462954 248294 463574 248378
rect 462954 248058 462986 248294
rect 463222 248058 463306 248294
rect 463542 248058 463574 248294
rect 462954 212614 463574 248058
rect 462954 212378 462986 212614
rect 463222 212378 463306 212614
rect 463542 212378 463574 212614
rect 462954 212294 463574 212378
rect 462954 212058 462986 212294
rect 463222 212058 463306 212294
rect 463542 212058 463574 212294
rect 462954 176614 463574 212058
rect 462954 176378 462986 176614
rect 463222 176378 463306 176614
rect 463542 176378 463574 176614
rect 462954 176294 463574 176378
rect 462954 176058 462986 176294
rect 463222 176058 463306 176294
rect 463542 176058 463574 176294
rect 462954 140614 463574 176058
rect 462954 140378 462986 140614
rect 463222 140378 463306 140614
rect 463542 140378 463574 140614
rect 462954 140294 463574 140378
rect 462954 140058 462986 140294
rect 463222 140058 463306 140294
rect 463542 140058 463574 140294
rect 462954 104614 463574 140058
rect 462954 104378 462986 104614
rect 463222 104378 463306 104614
rect 463542 104378 463574 104614
rect 462954 104294 463574 104378
rect 462954 104058 462986 104294
rect 463222 104058 463306 104294
rect 463542 104058 463574 104294
rect 462954 68614 463574 104058
rect 462954 68378 462986 68614
rect 463222 68378 463306 68614
rect 463542 68378 463574 68614
rect 462954 68294 463574 68378
rect 462954 68058 462986 68294
rect 463222 68058 463306 68294
rect 463542 68058 463574 68294
rect 462954 32614 463574 68058
rect 462954 32378 462986 32614
rect 463222 32378 463306 32614
rect 463542 32378 463574 32614
rect 462954 32294 463574 32378
rect 462954 32058 462986 32294
rect 463222 32058 463306 32294
rect 463542 32058 463574 32294
rect 444954 -6342 444986 -6106
rect 445222 -6342 445306 -6106
rect 445542 -6342 445574 -6106
rect 444954 -6426 445574 -6342
rect 444954 -6662 444986 -6426
rect 445222 -6662 445306 -6426
rect 445542 -6662 445574 -6426
rect 444954 -7654 445574 -6662
rect 462954 -7066 463574 32058
rect 469794 704838 470414 705830
rect 469794 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 470414 704838
rect 469794 704518 470414 704602
rect 469794 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 470414 704518
rect 469794 687454 470414 704282
rect 469794 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 470414 687454
rect 469794 687134 470414 687218
rect 469794 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 470414 687134
rect 469794 651454 470414 686898
rect 469794 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 470414 651454
rect 469794 651134 470414 651218
rect 469794 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 470414 651134
rect 469794 615454 470414 650898
rect 469794 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 470414 615454
rect 469794 615134 470414 615218
rect 469794 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 470414 615134
rect 469794 579454 470414 614898
rect 469794 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 470414 579454
rect 469794 579134 470414 579218
rect 469794 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 470414 579134
rect 469794 543454 470414 578898
rect 469794 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 470414 543454
rect 469794 543134 470414 543218
rect 469794 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 470414 543134
rect 469794 507454 470414 542898
rect 469794 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 470414 507454
rect 469794 507134 470414 507218
rect 469794 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 470414 507134
rect 469794 471454 470414 506898
rect 469794 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 470414 471454
rect 469794 471134 470414 471218
rect 469794 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 470414 471134
rect 469794 435454 470414 470898
rect 469794 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 470414 435454
rect 469794 435134 470414 435218
rect 469794 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 470414 435134
rect 469794 399454 470414 434898
rect 469794 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 470414 399454
rect 469794 399134 470414 399218
rect 469794 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 470414 399134
rect 469794 363454 470414 398898
rect 469794 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 470414 363454
rect 469794 363134 470414 363218
rect 469794 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 470414 363134
rect 469794 327454 470414 362898
rect 469794 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 470414 327454
rect 469794 327134 470414 327218
rect 469794 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 470414 327134
rect 469794 291454 470414 326898
rect 469794 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 470414 291454
rect 469794 291134 470414 291218
rect 469794 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 470414 291134
rect 469794 255454 470414 290898
rect 469794 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 470414 255454
rect 469794 255134 470414 255218
rect 469794 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 470414 255134
rect 469794 219454 470414 254898
rect 469794 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 470414 219454
rect 469794 219134 470414 219218
rect 469794 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 470414 219134
rect 469794 183454 470414 218898
rect 469794 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 470414 183454
rect 469794 183134 470414 183218
rect 469794 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 470414 183134
rect 469794 147454 470414 182898
rect 469794 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 470414 147454
rect 469794 147134 470414 147218
rect 469794 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 470414 147134
rect 469794 111454 470414 146898
rect 469794 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 470414 111454
rect 469794 111134 470414 111218
rect 469794 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 470414 111134
rect 469794 75454 470414 110898
rect 469794 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 470414 75454
rect 469794 75134 470414 75218
rect 469794 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 470414 75134
rect 469794 39454 470414 74898
rect 469794 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 470414 39454
rect 469794 39134 470414 39218
rect 469794 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 470414 39134
rect 469794 3454 470414 38898
rect 469794 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 470414 3454
rect 469794 3134 470414 3218
rect 469794 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 470414 3134
rect 469794 -346 470414 2898
rect 469794 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 470414 -346
rect 469794 -666 470414 -582
rect 469794 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 470414 -666
rect 469794 -1894 470414 -902
rect 473514 691174 474134 706202
rect 473514 690938 473546 691174
rect 473782 690938 473866 691174
rect 474102 690938 474134 691174
rect 473514 690854 474134 690938
rect 473514 690618 473546 690854
rect 473782 690618 473866 690854
rect 474102 690618 474134 690854
rect 473514 655174 474134 690618
rect 473514 654938 473546 655174
rect 473782 654938 473866 655174
rect 474102 654938 474134 655174
rect 473514 654854 474134 654938
rect 473514 654618 473546 654854
rect 473782 654618 473866 654854
rect 474102 654618 474134 654854
rect 473514 619174 474134 654618
rect 473514 618938 473546 619174
rect 473782 618938 473866 619174
rect 474102 618938 474134 619174
rect 473514 618854 474134 618938
rect 473514 618618 473546 618854
rect 473782 618618 473866 618854
rect 474102 618618 474134 618854
rect 473514 583174 474134 618618
rect 473514 582938 473546 583174
rect 473782 582938 473866 583174
rect 474102 582938 474134 583174
rect 473514 582854 474134 582938
rect 473514 582618 473546 582854
rect 473782 582618 473866 582854
rect 474102 582618 474134 582854
rect 473514 547174 474134 582618
rect 473514 546938 473546 547174
rect 473782 546938 473866 547174
rect 474102 546938 474134 547174
rect 473514 546854 474134 546938
rect 473514 546618 473546 546854
rect 473782 546618 473866 546854
rect 474102 546618 474134 546854
rect 473514 511174 474134 546618
rect 473514 510938 473546 511174
rect 473782 510938 473866 511174
rect 474102 510938 474134 511174
rect 473514 510854 474134 510938
rect 473514 510618 473546 510854
rect 473782 510618 473866 510854
rect 474102 510618 474134 510854
rect 473514 475174 474134 510618
rect 473514 474938 473546 475174
rect 473782 474938 473866 475174
rect 474102 474938 474134 475174
rect 473514 474854 474134 474938
rect 473514 474618 473546 474854
rect 473782 474618 473866 474854
rect 474102 474618 474134 474854
rect 473514 439174 474134 474618
rect 473514 438938 473546 439174
rect 473782 438938 473866 439174
rect 474102 438938 474134 439174
rect 473514 438854 474134 438938
rect 473514 438618 473546 438854
rect 473782 438618 473866 438854
rect 474102 438618 474134 438854
rect 473514 403174 474134 438618
rect 473514 402938 473546 403174
rect 473782 402938 473866 403174
rect 474102 402938 474134 403174
rect 473514 402854 474134 402938
rect 473514 402618 473546 402854
rect 473782 402618 473866 402854
rect 474102 402618 474134 402854
rect 473514 367174 474134 402618
rect 473514 366938 473546 367174
rect 473782 366938 473866 367174
rect 474102 366938 474134 367174
rect 473514 366854 474134 366938
rect 473514 366618 473546 366854
rect 473782 366618 473866 366854
rect 474102 366618 474134 366854
rect 473514 331174 474134 366618
rect 473514 330938 473546 331174
rect 473782 330938 473866 331174
rect 474102 330938 474134 331174
rect 473514 330854 474134 330938
rect 473514 330618 473546 330854
rect 473782 330618 473866 330854
rect 474102 330618 474134 330854
rect 473514 295174 474134 330618
rect 473514 294938 473546 295174
rect 473782 294938 473866 295174
rect 474102 294938 474134 295174
rect 473514 294854 474134 294938
rect 473514 294618 473546 294854
rect 473782 294618 473866 294854
rect 474102 294618 474134 294854
rect 473514 259174 474134 294618
rect 473514 258938 473546 259174
rect 473782 258938 473866 259174
rect 474102 258938 474134 259174
rect 473514 258854 474134 258938
rect 473514 258618 473546 258854
rect 473782 258618 473866 258854
rect 474102 258618 474134 258854
rect 473514 223174 474134 258618
rect 473514 222938 473546 223174
rect 473782 222938 473866 223174
rect 474102 222938 474134 223174
rect 473514 222854 474134 222938
rect 473514 222618 473546 222854
rect 473782 222618 473866 222854
rect 474102 222618 474134 222854
rect 473514 187174 474134 222618
rect 473514 186938 473546 187174
rect 473782 186938 473866 187174
rect 474102 186938 474134 187174
rect 473514 186854 474134 186938
rect 473514 186618 473546 186854
rect 473782 186618 473866 186854
rect 474102 186618 474134 186854
rect 473514 151174 474134 186618
rect 473514 150938 473546 151174
rect 473782 150938 473866 151174
rect 474102 150938 474134 151174
rect 473514 150854 474134 150938
rect 473514 150618 473546 150854
rect 473782 150618 473866 150854
rect 474102 150618 474134 150854
rect 473514 115174 474134 150618
rect 473514 114938 473546 115174
rect 473782 114938 473866 115174
rect 474102 114938 474134 115174
rect 473514 114854 474134 114938
rect 473514 114618 473546 114854
rect 473782 114618 473866 114854
rect 474102 114618 474134 114854
rect 473514 79174 474134 114618
rect 473514 78938 473546 79174
rect 473782 78938 473866 79174
rect 474102 78938 474134 79174
rect 473514 78854 474134 78938
rect 473514 78618 473546 78854
rect 473782 78618 473866 78854
rect 474102 78618 474134 78854
rect 473514 43174 474134 78618
rect 473514 42938 473546 43174
rect 473782 42938 473866 43174
rect 474102 42938 474134 43174
rect 473514 42854 474134 42938
rect 473514 42618 473546 42854
rect 473782 42618 473866 42854
rect 474102 42618 474134 42854
rect 473514 7174 474134 42618
rect 473514 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 474134 7174
rect 473514 6854 474134 6938
rect 473514 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 474134 6854
rect 473514 -2266 474134 6618
rect 473514 -2502 473546 -2266
rect 473782 -2502 473866 -2266
rect 474102 -2502 474134 -2266
rect 473514 -2586 474134 -2502
rect 473514 -2822 473546 -2586
rect 473782 -2822 473866 -2586
rect 474102 -2822 474134 -2586
rect 473514 -3814 474134 -2822
rect 477234 694894 477854 708122
rect 477234 694658 477266 694894
rect 477502 694658 477586 694894
rect 477822 694658 477854 694894
rect 477234 694574 477854 694658
rect 477234 694338 477266 694574
rect 477502 694338 477586 694574
rect 477822 694338 477854 694574
rect 477234 658894 477854 694338
rect 477234 658658 477266 658894
rect 477502 658658 477586 658894
rect 477822 658658 477854 658894
rect 477234 658574 477854 658658
rect 477234 658338 477266 658574
rect 477502 658338 477586 658574
rect 477822 658338 477854 658574
rect 477234 622894 477854 658338
rect 477234 622658 477266 622894
rect 477502 622658 477586 622894
rect 477822 622658 477854 622894
rect 477234 622574 477854 622658
rect 477234 622338 477266 622574
rect 477502 622338 477586 622574
rect 477822 622338 477854 622574
rect 477234 586894 477854 622338
rect 477234 586658 477266 586894
rect 477502 586658 477586 586894
rect 477822 586658 477854 586894
rect 477234 586574 477854 586658
rect 477234 586338 477266 586574
rect 477502 586338 477586 586574
rect 477822 586338 477854 586574
rect 477234 550894 477854 586338
rect 477234 550658 477266 550894
rect 477502 550658 477586 550894
rect 477822 550658 477854 550894
rect 477234 550574 477854 550658
rect 477234 550338 477266 550574
rect 477502 550338 477586 550574
rect 477822 550338 477854 550574
rect 477234 514894 477854 550338
rect 477234 514658 477266 514894
rect 477502 514658 477586 514894
rect 477822 514658 477854 514894
rect 477234 514574 477854 514658
rect 477234 514338 477266 514574
rect 477502 514338 477586 514574
rect 477822 514338 477854 514574
rect 477234 478894 477854 514338
rect 477234 478658 477266 478894
rect 477502 478658 477586 478894
rect 477822 478658 477854 478894
rect 477234 478574 477854 478658
rect 477234 478338 477266 478574
rect 477502 478338 477586 478574
rect 477822 478338 477854 478574
rect 477234 442894 477854 478338
rect 477234 442658 477266 442894
rect 477502 442658 477586 442894
rect 477822 442658 477854 442894
rect 477234 442574 477854 442658
rect 477234 442338 477266 442574
rect 477502 442338 477586 442574
rect 477822 442338 477854 442574
rect 477234 406894 477854 442338
rect 477234 406658 477266 406894
rect 477502 406658 477586 406894
rect 477822 406658 477854 406894
rect 477234 406574 477854 406658
rect 477234 406338 477266 406574
rect 477502 406338 477586 406574
rect 477822 406338 477854 406574
rect 477234 370894 477854 406338
rect 477234 370658 477266 370894
rect 477502 370658 477586 370894
rect 477822 370658 477854 370894
rect 477234 370574 477854 370658
rect 477234 370338 477266 370574
rect 477502 370338 477586 370574
rect 477822 370338 477854 370574
rect 477234 334894 477854 370338
rect 477234 334658 477266 334894
rect 477502 334658 477586 334894
rect 477822 334658 477854 334894
rect 477234 334574 477854 334658
rect 477234 334338 477266 334574
rect 477502 334338 477586 334574
rect 477822 334338 477854 334574
rect 477234 298894 477854 334338
rect 477234 298658 477266 298894
rect 477502 298658 477586 298894
rect 477822 298658 477854 298894
rect 477234 298574 477854 298658
rect 477234 298338 477266 298574
rect 477502 298338 477586 298574
rect 477822 298338 477854 298574
rect 477234 262894 477854 298338
rect 477234 262658 477266 262894
rect 477502 262658 477586 262894
rect 477822 262658 477854 262894
rect 477234 262574 477854 262658
rect 477234 262338 477266 262574
rect 477502 262338 477586 262574
rect 477822 262338 477854 262574
rect 477234 226894 477854 262338
rect 477234 226658 477266 226894
rect 477502 226658 477586 226894
rect 477822 226658 477854 226894
rect 477234 226574 477854 226658
rect 477234 226338 477266 226574
rect 477502 226338 477586 226574
rect 477822 226338 477854 226574
rect 477234 190894 477854 226338
rect 477234 190658 477266 190894
rect 477502 190658 477586 190894
rect 477822 190658 477854 190894
rect 477234 190574 477854 190658
rect 477234 190338 477266 190574
rect 477502 190338 477586 190574
rect 477822 190338 477854 190574
rect 477234 154894 477854 190338
rect 477234 154658 477266 154894
rect 477502 154658 477586 154894
rect 477822 154658 477854 154894
rect 477234 154574 477854 154658
rect 477234 154338 477266 154574
rect 477502 154338 477586 154574
rect 477822 154338 477854 154574
rect 477234 118894 477854 154338
rect 477234 118658 477266 118894
rect 477502 118658 477586 118894
rect 477822 118658 477854 118894
rect 477234 118574 477854 118658
rect 477234 118338 477266 118574
rect 477502 118338 477586 118574
rect 477822 118338 477854 118574
rect 477234 82894 477854 118338
rect 477234 82658 477266 82894
rect 477502 82658 477586 82894
rect 477822 82658 477854 82894
rect 477234 82574 477854 82658
rect 477234 82338 477266 82574
rect 477502 82338 477586 82574
rect 477822 82338 477854 82574
rect 477234 46894 477854 82338
rect 477234 46658 477266 46894
rect 477502 46658 477586 46894
rect 477822 46658 477854 46894
rect 477234 46574 477854 46658
rect 477234 46338 477266 46574
rect 477502 46338 477586 46574
rect 477822 46338 477854 46574
rect 477234 10894 477854 46338
rect 477234 10658 477266 10894
rect 477502 10658 477586 10894
rect 477822 10658 477854 10894
rect 477234 10574 477854 10658
rect 477234 10338 477266 10574
rect 477502 10338 477586 10574
rect 477822 10338 477854 10574
rect 477234 -4186 477854 10338
rect 477234 -4422 477266 -4186
rect 477502 -4422 477586 -4186
rect 477822 -4422 477854 -4186
rect 477234 -4506 477854 -4422
rect 477234 -4742 477266 -4506
rect 477502 -4742 477586 -4506
rect 477822 -4742 477854 -4506
rect 477234 -5734 477854 -4742
rect 480954 698614 481574 710042
rect 498954 711558 499574 711590
rect 498954 711322 498986 711558
rect 499222 711322 499306 711558
rect 499542 711322 499574 711558
rect 498954 711238 499574 711322
rect 498954 711002 498986 711238
rect 499222 711002 499306 711238
rect 499542 711002 499574 711238
rect 495234 709638 495854 709670
rect 495234 709402 495266 709638
rect 495502 709402 495586 709638
rect 495822 709402 495854 709638
rect 495234 709318 495854 709402
rect 495234 709082 495266 709318
rect 495502 709082 495586 709318
rect 495822 709082 495854 709318
rect 491514 707718 492134 707750
rect 491514 707482 491546 707718
rect 491782 707482 491866 707718
rect 492102 707482 492134 707718
rect 491514 707398 492134 707482
rect 491514 707162 491546 707398
rect 491782 707162 491866 707398
rect 492102 707162 492134 707398
rect 480954 698378 480986 698614
rect 481222 698378 481306 698614
rect 481542 698378 481574 698614
rect 480954 698294 481574 698378
rect 480954 698058 480986 698294
rect 481222 698058 481306 698294
rect 481542 698058 481574 698294
rect 480954 662614 481574 698058
rect 480954 662378 480986 662614
rect 481222 662378 481306 662614
rect 481542 662378 481574 662614
rect 480954 662294 481574 662378
rect 480954 662058 480986 662294
rect 481222 662058 481306 662294
rect 481542 662058 481574 662294
rect 480954 626614 481574 662058
rect 480954 626378 480986 626614
rect 481222 626378 481306 626614
rect 481542 626378 481574 626614
rect 480954 626294 481574 626378
rect 480954 626058 480986 626294
rect 481222 626058 481306 626294
rect 481542 626058 481574 626294
rect 480954 590614 481574 626058
rect 480954 590378 480986 590614
rect 481222 590378 481306 590614
rect 481542 590378 481574 590614
rect 480954 590294 481574 590378
rect 480954 590058 480986 590294
rect 481222 590058 481306 590294
rect 481542 590058 481574 590294
rect 480954 554614 481574 590058
rect 480954 554378 480986 554614
rect 481222 554378 481306 554614
rect 481542 554378 481574 554614
rect 480954 554294 481574 554378
rect 480954 554058 480986 554294
rect 481222 554058 481306 554294
rect 481542 554058 481574 554294
rect 480954 518614 481574 554058
rect 480954 518378 480986 518614
rect 481222 518378 481306 518614
rect 481542 518378 481574 518614
rect 480954 518294 481574 518378
rect 480954 518058 480986 518294
rect 481222 518058 481306 518294
rect 481542 518058 481574 518294
rect 480954 482614 481574 518058
rect 480954 482378 480986 482614
rect 481222 482378 481306 482614
rect 481542 482378 481574 482614
rect 480954 482294 481574 482378
rect 480954 482058 480986 482294
rect 481222 482058 481306 482294
rect 481542 482058 481574 482294
rect 480954 446614 481574 482058
rect 480954 446378 480986 446614
rect 481222 446378 481306 446614
rect 481542 446378 481574 446614
rect 480954 446294 481574 446378
rect 480954 446058 480986 446294
rect 481222 446058 481306 446294
rect 481542 446058 481574 446294
rect 480954 410614 481574 446058
rect 480954 410378 480986 410614
rect 481222 410378 481306 410614
rect 481542 410378 481574 410614
rect 480954 410294 481574 410378
rect 480954 410058 480986 410294
rect 481222 410058 481306 410294
rect 481542 410058 481574 410294
rect 480954 374614 481574 410058
rect 480954 374378 480986 374614
rect 481222 374378 481306 374614
rect 481542 374378 481574 374614
rect 480954 374294 481574 374378
rect 480954 374058 480986 374294
rect 481222 374058 481306 374294
rect 481542 374058 481574 374294
rect 480954 338614 481574 374058
rect 480954 338378 480986 338614
rect 481222 338378 481306 338614
rect 481542 338378 481574 338614
rect 480954 338294 481574 338378
rect 480954 338058 480986 338294
rect 481222 338058 481306 338294
rect 481542 338058 481574 338294
rect 480954 302614 481574 338058
rect 480954 302378 480986 302614
rect 481222 302378 481306 302614
rect 481542 302378 481574 302614
rect 480954 302294 481574 302378
rect 480954 302058 480986 302294
rect 481222 302058 481306 302294
rect 481542 302058 481574 302294
rect 480954 266614 481574 302058
rect 480954 266378 480986 266614
rect 481222 266378 481306 266614
rect 481542 266378 481574 266614
rect 480954 266294 481574 266378
rect 480954 266058 480986 266294
rect 481222 266058 481306 266294
rect 481542 266058 481574 266294
rect 480954 230614 481574 266058
rect 480954 230378 480986 230614
rect 481222 230378 481306 230614
rect 481542 230378 481574 230614
rect 480954 230294 481574 230378
rect 480954 230058 480986 230294
rect 481222 230058 481306 230294
rect 481542 230058 481574 230294
rect 480954 194614 481574 230058
rect 480954 194378 480986 194614
rect 481222 194378 481306 194614
rect 481542 194378 481574 194614
rect 480954 194294 481574 194378
rect 480954 194058 480986 194294
rect 481222 194058 481306 194294
rect 481542 194058 481574 194294
rect 480954 158614 481574 194058
rect 480954 158378 480986 158614
rect 481222 158378 481306 158614
rect 481542 158378 481574 158614
rect 480954 158294 481574 158378
rect 480954 158058 480986 158294
rect 481222 158058 481306 158294
rect 481542 158058 481574 158294
rect 480954 122614 481574 158058
rect 480954 122378 480986 122614
rect 481222 122378 481306 122614
rect 481542 122378 481574 122614
rect 480954 122294 481574 122378
rect 480954 122058 480986 122294
rect 481222 122058 481306 122294
rect 481542 122058 481574 122294
rect 480954 86614 481574 122058
rect 480954 86378 480986 86614
rect 481222 86378 481306 86614
rect 481542 86378 481574 86614
rect 480954 86294 481574 86378
rect 480954 86058 480986 86294
rect 481222 86058 481306 86294
rect 481542 86058 481574 86294
rect 480954 50614 481574 86058
rect 480954 50378 480986 50614
rect 481222 50378 481306 50614
rect 481542 50378 481574 50614
rect 480954 50294 481574 50378
rect 480954 50058 480986 50294
rect 481222 50058 481306 50294
rect 481542 50058 481574 50294
rect 480954 14614 481574 50058
rect 480954 14378 480986 14614
rect 481222 14378 481306 14614
rect 481542 14378 481574 14614
rect 480954 14294 481574 14378
rect 480954 14058 480986 14294
rect 481222 14058 481306 14294
rect 481542 14058 481574 14294
rect 462954 -7302 462986 -7066
rect 463222 -7302 463306 -7066
rect 463542 -7302 463574 -7066
rect 462954 -7386 463574 -7302
rect 462954 -7622 462986 -7386
rect 463222 -7622 463306 -7386
rect 463542 -7622 463574 -7386
rect 462954 -7654 463574 -7622
rect 480954 -6106 481574 14058
rect 487794 705798 488414 705830
rect 487794 705562 487826 705798
rect 488062 705562 488146 705798
rect 488382 705562 488414 705798
rect 487794 705478 488414 705562
rect 487794 705242 487826 705478
rect 488062 705242 488146 705478
rect 488382 705242 488414 705478
rect 487794 669454 488414 705242
rect 487794 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 488414 669454
rect 487794 669134 488414 669218
rect 487794 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 488414 669134
rect 487794 633454 488414 668898
rect 487794 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 488414 633454
rect 487794 633134 488414 633218
rect 487794 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 488414 633134
rect 487794 597454 488414 632898
rect 487794 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 488414 597454
rect 487794 597134 488414 597218
rect 487794 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 488414 597134
rect 487794 561454 488414 596898
rect 487794 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 488414 561454
rect 487794 561134 488414 561218
rect 487794 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 488414 561134
rect 487794 525454 488414 560898
rect 487794 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 488414 525454
rect 487794 525134 488414 525218
rect 487794 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 488414 525134
rect 487794 489454 488414 524898
rect 487794 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 488414 489454
rect 487794 489134 488414 489218
rect 487794 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 488414 489134
rect 487794 453454 488414 488898
rect 487794 453218 487826 453454
rect 488062 453218 488146 453454
rect 488382 453218 488414 453454
rect 487794 453134 488414 453218
rect 487794 452898 487826 453134
rect 488062 452898 488146 453134
rect 488382 452898 488414 453134
rect 487794 417454 488414 452898
rect 487794 417218 487826 417454
rect 488062 417218 488146 417454
rect 488382 417218 488414 417454
rect 487794 417134 488414 417218
rect 487794 416898 487826 417134
rect 488062 416898 488146 417134
rect 488382 416898 488414 417134
rect 487794 381454 488414 416898
rect 487794 381218 487826 381454
rect 488062 381218 488146 381454
rect 488382 381218 488414 381454
rect 487794 381134 488414 381218
rect 487794 380898 487826 381134
rect 488062 380898 488146 381134
rect 488382 380898 488414 381134
rect 487794 345454 488414 380898
rect 487794 345218 487826 345454
rect 488062 345218 488146 345454
rect 488382 345218 488414 345454
rect 487794 345134 488414 345218
rect 487794 344898 487826 345134
rect 488062 344898 488146 345134
rect 488382 344898 488414 345134
rect 487794 309454 488414 344898
rect 487794 309218 487826 309454
rect 488062 309218 488146 309454
rect 488382 309218 488414 309454
rect 487794 309134 488414 309218
rect 487794 308898 487826 309134
rect 488062 308898 488146 309134
rect 488382 308898 488414 309134
rect 487794 273454 488414 308898
rect 487794 273218 487826 273454
rect 488062 273218 488146 273454
rect 488382 273218 488414 273454
rect 487794 273134 488414 273218
rect 487794 272898 487826 273134
rect 488062 272898 488146 273134
rect 488382 272898 488414 273134
rect 487794 237454 488414 272898
rect 487794 237218 487826 237454
rect 488062 237218 488146 237454
rect 488382 237218 488414 237454
rect 487794 237134 488414 237218
rect 487794 236898 487826 237134
rect 488062 236898 488146 237134
rect 488382 236898 488414 237134
rect 487794 201454 488414 236898
rect 487794 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 488414 201454
rect 487794 201134 488414 201218
rect 487794 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 488414 201134
rect 487794 165454 488414 200898
rect 487794 165218 487826 165454
rect 488062 165218 488146 165454
rect 488382 165218 488414 165454
rect 487794 165134 488414 165218
rect 487794 164898 487826 165134
rect 488062 164898 488146 165134
rect 488382 164898 488414 165134
rect 487794 129454 488414 164898
rect 487794 129218 487826 129454
rect 488062 129218 488146 129454
rect 488382 129218 488414 129454
rect 487794 129134 488414 129218
rect 487794 128898 487826 129134
rect 488062 128898 488146 129134
rect 488382 128898 488414 129134
rect 487794 93454 488414 128898
rect 487794 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 488414 93454
rect 487794 93134 488414 93218
rect 487794 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 488414 93134
rect 487794 57454 488414 92898
rect 487794 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 488414 57454
rect 487794 57134 488414 57218
rect 487794 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 488414 57134
rect 487794 21454 488414 56898
rect 487794 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 488414 21454
rect 487794 21134 488414 21218
rect 487794 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 488414 21134
rect 487794 -1306 488414 20898
rect 487794 -1542 487826 -1306
rect 488062 -1542 488146 -1306
rect 488382 -1542 488414 -1306
rect 487794 -1626 488414 -1542
rect 487794 -1862 487826 -1626
rect 488062 -1862 488146 -1626
rect 488382 -1862 488414 -1626
rect 487794 -1894 488414 -1862
rect 491514 673174 492134 707162
rect 491514 672938 491546 673174
rect 491782 672938 491866 673174
rect 492102 672938 492134 673174
rect 491514 672854 492134 672938
rect 491514 672618 491546 672854
rect 491782 672618 491866 672854
rect 492102 672618 492134 672854
rect 491514 637174 492134 672618
rect 491514 636938 491546 637174
rect 491782 636938 491866 637174
rect 492102 636938 492134 637174
rect 491514 636854 492134 636938
rect 491514 636618 491546 636854
rect 491782 636618 491866 636854
rect 492102 636618 492134 636854
rect 491514 601174 492134 636618
rect 491514 600938 491546 601174
rect 491782 600938 491866 601174
rect 492102 600938 492134 601174
rect 491514 600854 492134 600938
rect 491514 600618 491546 600854
rect 491782 600618 491866 600854
rect 492102 600618 492134 600854
rect 491514 565174 492134 600618
rect 491514 564938 491546 565174
rect 491782 564938 491866 565174
rect 492102 564938 492134 565174
rect 491514 564854 492134 564938
rect 491514 564618 491546 564854
rect 491782 564618 491866 564854
rect 492102 564618 492134 564854
rect 491514 529174 492134 564618
rect 491514 528938 491546 529174
rect 491782 528938 491866 529174
rect 492102 528938 492134 529174
rect 491514 528854 492134 528938
rect 491514 528618 491546 528854
rect 491782 528618 491866 528854
rect 492102 528618 492134 528854
rect 491514 493174 492134 528618
rect 491514 492938 491546 493174
rect 491782 492938 491866 493174
rect 492102 492938 492134 493174
rect 491514 492854 492134 492938
rect 491514 492618 491546 492854
rect 491782 492618 491866 492854
rect 492102 492618 492134 492854
rect 491514 457174 492134 492618
rect 491514 456938 491546 457174
rect 491782 456938 491866 457174
rect 492102 456938 492134 457174
rect 491514 456854 492134 456938
rect 491514 456618 491546 456854
rect 491782 456618 491866 456854
rect 492102 456618 492134 456854
rect 491514 421174 492134 456618
rect 491514 420938 491546 421174
rect 491782 420938 491866 421174
rect 492102 420938 492134 421174
rect 491514 420854 492134 420938
rect 491514 420618 491546 420854
rect 491782 420618 491866 420854
rect 492102 420618 492134 420854
rect 491514 385174 492134 420618
rect 491514 384938 491546 385174
rect 491782 384938 491866 385174
rect 492102 384938 492134 385174
rect 491514 384854 492134 384938
rect 491514 384618 491546 384854
rect 491782 384618 491866 384854
rect 492102 384618 492134 384854
rect 491514 349174 492134 384618
rect 491514 348938 491546 349174
rect 491782 348938 491866 349174
rect 492102 348938 492134 349174
rect 491514 348854 492134 348938
rect 491514 348618 491546 348854
rect 491782 348618 491866 348854
rect 492102 348618 492134 348854
rect 491514 313174 492134 348618
rect 491514 312938 491546 313174
rect 491782 312938 491866 313174
rect 492102 312938 492134 313174
rect 491514 312854 492134 312938
rect 491514 312618 491546 312854
rect 491782 312618 491866 312854
rect 492102 312618 492134 312854
rect 491514 277174 492134 312618
rect 491514 276938 491546 277174
rect 491782 276938 491866 277174
rect 492102 276938 492134 277174
rect 491514 276854 492134 276938
rect 491514 276618 491546 276854
rect 491782 276618 491866 276854
rect 492102 276618 492134 276854
rect 491514 241174 492134 276618
rect 491514 240938 491546 241174
rect 491782 240938 491866 241174
rect 492102 240938 492134 241174
rect 491514 240854 492134 240938
rect 491514 240618 491546 240854
rect 491782 240618 491866 240854
rect 492102 240618 492134 240854
rect 491514 205174 492134 240618
rect 491514 204938 491546 205174
rect 491782 204938 491866 205174
rect 492102 204938 492134 205174
rect 491514 204854 492134 204938
rect 491514 204618 491546 204854
rect 491782 204618 491866 204854
rect 492102 204618 492134 204854
rect 491514 169174 492134 204618
rect 491514 168938 491546 169174
rect 491782 168938 491866 169174
rect 492102 168938 492134 169174
rect 491514 168854 492134 168938
rect 491514 168618 491546 168854
rect 491782 168618 491866 168854
rect 492102 168618 492134 168854
rect 491514 133174 492134 168618
rect 491514 132938 491546 133174
rect 491782 132938 491866 133174
rect 492102 132938 492134 133174
rect 491514 132854 492134 132938
rect 491514 132618 491546 132854
rect 491782 132618 491866 132854
rect 492102 132618 492134 132854
rect 491514 97174 492134 132618
rect 491514 96938 491546 97174
rect 491782 96938 491866 97174
rect 492102 96938 492134 97174
rect 491514 96854 492134 96938
rect 491514 96618 491546 96854
rect 491782 96618 491866 96854
rect 492102 96618 492134 96854
rect 491514 61174 492134 96618
rect 491514 60938 491546 61174
rect 491782 60938 491866 61174
rect 492102 60938 492134 61174
rect 491514 60854 492134 60938
rect 491514 60618 491546 60854
rect 491782 60618 491866 60854
rect 492102 60618 492134 60854
rect 491514 25174 492134 60618
rect 491514 24938 491546 25174
rect 491782 24938 491866 25174
rect 492102 24938 492134 25174
rect 491514 24854 492134 24938
rect 491514 24618 491546 24854
rect 491782 24618 491866 24854
rect 492102 24618 492134 24854
rect 491514 -3226 492134 24618
rect 491514 -3462 491546 -3226
rect 491782 -3462 491866 -3226
rect 492102 -3462 492134 -3226
rect 491514 -3546 492134 -3462
rect 491514 -3782 491546 -3546
rect 491782 -3782 491866 -3546
rect 492102 -3782 492134 -3546
rect 491514 -3814 492134 -3782
rect 495234 676894 495854 709082
rect 495234 676658 495266 676894
rect 495502 676658 495586 676894
rect 495822 676658 495854 676894
rect 495234 676574 495854 676658
rect 495234 676338 495266 676574
rect 495502 676338 495586 676574
rect 495822 676338 495854 676574
rect 495234 640894 495854 676338
rect 495234 640658 495266 640894
rect 495502 640658 495586 640894
rect 495822 640658 495854 640894
rect 495234 640574 495854 640658
rect 495234 640338 495266 640574
rect 495502 640338 495586 640574
rect 495822 640338 495854 640574
rect 495234 604894 495854 640338
rect 495234 604658 495266 604894
rect 495502 604658 495586 604894
rect 495822 604658 495854 604894
rect 495234 604574 495854 604658
rect 495234 604338 495266 604574
rect 495502 604338 495586 604574
rect 495822 604338 495854 604574
rect 495234 568894 495854 604338
rect 495234 568658 495266 568894
rect 495502 568658 495586 568894
rect 495822 568658 495854 568894
rect 495234 568574 495854 568658
rect 495234 568338 495266 568574
rect 495502 568338 495586 568574
rect 495822 568338 495854 568574
rect 495234 532894 495854 568338
rect 495234 532658 495266 532894
rect 495502 532658 495586 532894
rect 495822 532658 495854 532894
rect 495234 532574 495854 532658
rect 495234 532338 495266 532574
rect 495502 532338 495586 532574
rect 495822 532338 495854 532574
rect 495234 496894 495854 532338
rect 495234 496658 495266 496894
rect 495502 496658 495586 496894
rect 495822 496658 495854 496894
rect 495234 496574 495854 496658
rect 495234 496338 495266 496574
rect 495502 496338 495586 496574
rect 495822 496338 495854 496574
rect 495234 460894 495854 496338
rect 495234 460658 495266 460894
rect 495502 460658 495586 460894
rect 495822 460658 495854 460894
rect 495234 460574 495854 460658
rect 495234 460338 495266 460574
rect 495502 460338 495586 460574
rect 495822 460338 495854 460574
rect 495234 424894 495854 460338
rect 495234 424658 495266 424894
rect 495502 424658 495586 424894
rect 495822 424658 495854 424894
rect 495234 424574 495854 424658
rect 495234 424338 495266 424574
rect 495502 424338 495586 424574
rect 495822 424338 495854 424574
rect 495234 388894 495854 424338
rect 495234 388658 495266 388894
rect 495502 388658 495586 388894
rect 495822 388658 495854 388894
rect 495234 388574 495854 388658
rect 495234 388338 495266 388574
rect 495502 388338 495586 388574
rect 495822 388338 495854 388574
rect 495234 352894 495854 388338
rect 495234 352658 495266 352894
rect 495502 352658 495586 352894
rect 495822 352658 495854 352894
rect 495234 352574 495854 352658
rect 495234 352338 495266 352574
rect 495502 352338 495586 352574
rect 495822 352338 495854 352574
rect 495234 316894 495854 352338
rect 495234 316658 495266 316894
rect 495502 316658 495586 316894
rect 495822 316658 495854 316894
rect 495234 316574 495854 316658
rect 495234 316338 495266 316574
rect 495502 316338 495586 316574
rect 495822 316338 495854 316574
rect 495234 280894 495854 316338
rect 495234 280658 495266 280894
rect 495502 280658 495586 280894
rect 495822 280658 495854 280894
rect 495234 280574 495854 280658
rect 495234 280338 495266 280574
rect 495502 280338 495586 280574
rect 495822 280338 495854 280574
rect 495234 244894 495854 280338
rect 495234 244658 495266 244894
rect 495502 244658 495586 244894
rect 495822 244658 495854 244894
rect 495234 244574 495854 244658
rect 495234 244338 495266 244574
rect 495502 244338 495586 244574
rect 495822 244338 495854 244574
rect 495234 208894 495854 244338
rect 495234 208658 495266 208894
rect 495502 208658 495586 208894
rect 495822 208658 495854 208894
rect 495234 208574 495854 208658
rect 495234 208338 495266 208574
rect 495502 208338 495586 208574
rect 495822 208338 495854 208574
rect 495234 172894 495854 208338
rect 495234 172658 495266 172894
rect 495502 172658 495586 172894
rect 495822 172658 495854 172894
rect 495234 172574 495854 172658
rect 495234 172338 495266 172574
rect 495502 172338 495586 172574
rect 495822 172338 495854 172574
rect 495234 136894 495854 172338
rect 495234 136658 495266 136894
rect 495502 136658 495586 136894
rect 495822 136658 495854 136894
rect 495234 136574 495854 136658
rect 495234 136338 495266 136574
rect 495502 136338 495586 136574
rect 495822 136338 495854 136574
rect 495234 100894 495854 136338
rect 495234 100658 495266 100894
rect 495502 100658 495586 100894
rect 495822 100658 495854 100894
rect 495234 100574 495854 100658
rect 495234 100338 495266 100574
rect 495502 100338 495586 100574
rect 495822 100338 495854 100574
rect 495234 64894 495854 100338
rect 495234 64658 495266 64894
rect 495502 64658 495586 64894
rect 495822 64658 495854 64894
rect 495234 64574 495854 64658
rect 495234 64338 495266 64574
rect 495502 64338 495586 64574
rect 495822 64338 495854 64574
rect 495234 28894 495854 64338
rect 495234 28658 495266 28894
rect 495502 28658 495586 28894
rect 495822 28658 495854 28894
rect 495234 28574 495854 28658
rect 495234 28338 495266 28574
rect 495502 28338 495586 28574
rect 495822 28338 495854 28574
rect 495234 -5146 495854 28338
rect 495234 -5382 495266 -5146
rect 495502 -5382 495586 -5146
rect 495822 -5382 495854 -5146
rect 495234 -5466 495854 -5382
rect 495234 -5702 495266 -5466
rect 495502 -5702 495586 -5466
rect 495822 -5702 495854 -5466
rect 495234 -5734 495854 -5702
rect 498954 680614 499574 711002
rect 516954 710598 517574 711590
rect 516954 710362 516986 710598
rect 517222 710362 517306 710598
rect 517542 710362 517574 710598
rect 516954 710278 517574 710362
rect 516954 710042 516986 710278
rect 517222 710042 517306 710278
rect 517542 710042 517574 710278
rect 513234 708678 513854 709670
rect 513234 708442 513266 708678
rect 513502 708442 513586 708678
rect 513822 708442 513854 708678
rect 513234 708358 513854 708442
rect 513234 708122 513266 708358
rect 513502 708122 513586 708358
rect 513822 708122 513854 708358
rect 509514 706758 510134 707750
rect 509514 706522 509546 706758
rect 509782 706522 509866 706758
rect 510102 706522 510134 706758
rect 509514 706438 510134 706522
rect 509514 706202 509546 706438
rect 509782 706202 509866 706438
rect 510102 706202 510134 706438
rect 498954 680378 498986 680614
rect 499222 680378 499306 680614
rect 499542 680378 499574 680614
rect 498954 680294 499574 680378
rect 498954 680058 498986 680294
rect 499222 680058 499306 680294
rect 499542 680058 499574 680294
rect 498954 644614 499574 680058
rect 498954 644378 498986 644614
rect 499222 644378 499306 644614
rect 499542 644378 499574 644614
rect 498954 644294 499574 644378
rect 498954 644058 498986 644294
rect 499222 644058 499306 644294
rect 499542 644058 499574 644294
rect 498954 608614 499574 644058
rect 498954 608378 498986 608614
rect 499222 608378 499306 608614
rect 499542 608378 499574 608614
rect 498954 608294 499574 608378
rect 498954 608058 498986 608294
rect 499222 608058 499306 608294
rect 499542 608058 499574 608294
rect 498954 572614 499574 608058
rect 498954 572378 498986 572614
rect 499222 572378 499306 572614
rect 499542 572378 499574 572614
rect 498954 572294 499574 572378
rect 498954 572058 498986 572294
rect 499222 572058 499306 572294
rect 499542 572058 499574 572294
rect 498954 536614 499574 572058
rect 498954 536378 498986 536614
rect 499222 536378 499306 536614
rect 499542 536378 499574 536614
rect 498954 536294 499574 536378
rect 498954 536058 498986 536294
rect 499222 536058 499306 536294
rect 499542 536058 499574 536294
rect 498954 500614 499574 536058
rect 498954 500378 498986 500614
rect 499222 500378 499306 500614
rect 499542 500378 499574 500614
rect 498954 500294 499574 500378
rect 498954 500058 498986 500294
rect 499222 500058 499306 500294
rect 499542 500058 499574 500294
rect 498954 464614 499574 500058
rect 498954 464378 498986 464614
rect 499222 464378 499306 464614
rect 499542 464378 499574 464614
rect 498954 464294 499574 464378
rect 498954 464058 498986 464294
rect 499222 464058 499306 464294
rect 499542 464058 499574 464294
rect 498954 428614 499574 464058
rect 498954 428378 498986 428614
rect 499222 428378 499306 428614
rect 499542 428378 499574 428614
rect 498954 428294 499574 428378
rect 498954 428058 498986 428294
rect 499222 428058 499306 428294
rect 499542 428058 499574 428294
rect 498954 392614 499574 428058
rect 498954 392378 498986 392614
rect 499222 392378 499306 392614
rect 499542 392378 499574 392614
rect 498954 392294 499574 392378
rect 498954 392058 498986 392294
rect 499222 392058 499306 392294
rect 499542 392058 499574 392294
rect 498954 356614 499574 392058
rect 498954 356378 498986 356614
rect 499222 356378 499306 356614
rect 499542 356378 499574 356614
rect 498954 356294 499574 356378
rect 498954 356058 498986 356294
rect 499222 356058 499306 356294
rect 499542 356058 499574 356294
rect 498954 320614 499574 356058
rect 498954 320378 498986 320614
rect 499222 320378 499306 320614
rect 499542 320378 499574 320614
rect 498954 320294 499574 320378
rect 498954 320058 498986 320294
rect 499222 320058 499306 320294
rect 499542 320058 499574 320294
rect 498954 284614 499574 320058
rect 498954 284378 498986 284614
rect 499222 284378 499306 284614
rect 499542 284378 499574 284614
rect 498954 284294 499574 284378
rect 498954 284058 498986 284294
rect 499222 284058 499306 284294
rect 499542 284058 499574 284294
rect 498954 248614 499574 284058
rect 498954 248378 498986 248614
rect 499222 248378 499306 248614
rect 499542 248378 499574 248614
rect 498954 248294 499574 248378
rect 498954 248058 498986 248294
rect 499222 248058 499306 248294
rect 499542 248058 499574 248294
rect 498954 212614 499574 248058
rect 498954 212378 498986 212614
rect 499222 212378 499306 212614
rect 499542 212378 499574 212614
rect 498954 212294 499574 212378
rect 498954 212058 498986 212294
rect 499222 212058 499306 212294
rect 499542 212058 499574 212294
rect 498954 176614 499574 212058
rect 498954 176378 498986 176614
rect 499222 176378 499306 176614
rect 499542 176378 499574 176614
rect 498954 176294 499574 176378
rect 498954 176058 498986 176294
rect 499222 176058 499306 176294
rect 499542 176058 499574 176294
rect 498954 140614 499574 176058
rect 498954 140378 498986 140614
rect 499222 140378 499306 140614
rect 499542 140378 499574 140614
rect 498954 140294 499574 140378
rect 498954 140058 498986 140294
rect 499222 140058 499306 140294
rect 499542 140058 499574 140294
rect 498954 104614 499574 140058
rect 498954 104378 498986 104614
rect 499222 104378 499306 104614
rect 499542 104378 499574 104614
rect 498954 104294 499574 104378
rect 498954 104058 498986 104294
rect 499222 104058 499306 104294
rect 499542 104058 499574 104294
rect 498954 68614 499574 104058
rect 498954 68378 498986 68614
rect 499222 68378 499306 68614
rect 499542 68378 499574 68614
rect 498954 68294 499574 68378
rect 498954 68058 498986 68294
rect 499222 68058 499306 68294
rect 499542 68058 499574 68294
rect 498954 32614 499574 68058
rect 498954 32378 498986 32614
rect 499222 32378 499306 32614
rect 499542 32378 499574 32614
rect 498954 32294 499574 32378
rect 498954 32058 498986 32294
rect 499222 32058 499306 32294
rect 499542 32058 499574 32294
rect 480954 -6342 480986 -6106
rect 481222 -6342 481306 -6106
rect 481542 -6342 481574 -6106
rect 480954 -6426 481574 -6342
rect 480954 -6662 480986 -6426
rect 481222 -6662 481306 -6426
rect 481542 -6662 481574 -6426
rect 480954 -7654 481574 -6662
rect 498954 -7066 499574 32058
rect 505794 704838 506414 705830
rect 505794 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 506414 704838
rect 505794 704518 506414 704602
rect 505794 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 506414 704518
rect 505794 687454 506414 704282
rect 505794 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 506414 687454
rect 505794 687134 506414 687218
rect 505794 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 506414 687134
rect 505794 651454 506414 686898
rect 505794 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 506414 651454
rect 505794 651134 506414 651218
rect 505794 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 506414 651134
rect 505794 615454 506414 650898
rect 505794 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 506414 615454
rect 505794 615134 506414 615218
rect 505794 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 506414 615134
rect 505794 579454 506414 614898
rect 505794 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 506414 579454
rect 505794 579134 506414 579218
rect 505794 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 506414 579134
rect 505794 543454 506414 578898
rect 505794 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 506414 543454
rect 505794 543134 506414 543218
rect 505794 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 506414 543134
rect 505794 507454 506414 542898
rect 505794 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 506414 507454
rect 505794 507134 506414 507218
rect 505794 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 506414 507134
rect 505794 471454 506414 506898
rect 505794 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 506414 471454
rect 505794 471134 506414 471218
rect 505794 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 506414 471134
rect 505794 435454 506414 470898
rect 505794 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 506414 435454
rect 505794 435134 506414 435218
rect 505794 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 506414 435134
rect 505794 399454 506414 434898
rect 505794 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 506414 399454
rect 505794 399134 506414 399218
rect 505794 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 506414 399134
rect 505794 363454 506414 398898
rect 505794 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 506414 363454
rect 505794 363134 506414 363218
rect 505794 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 506414 363134
rect 505794 327454 506414 362898
rect 505794 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 506414 327454
rect 505794 327134 506414 327218
rect 505794 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 506414 327134
rect 505794 291454 506414 326898
rect 505794 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 506414 291454
rect 505794 291134 506414 291218
rect 505794 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 506414 291134
rect 505794 255454 506414 290898
rect 505794 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 506414 255454
rect 505794 255134 506414 255218
rect 505794 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 506414 255134
rect 505794 219454 506414 254898
rect 505794 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 506414 219454
rect 505794 219134 506414 219218
rect 505794 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 506414 219134
rect 505794 183454 506414 218898
rect 505794 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 506414 183454
rect 505794 183134 506414 183218
rect 505794 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 506414 183134
rect 505794 147454 506414 182898
rect 505794 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 506414 147454
rect 505794 147134 506414 147218
rect 505794 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 506414 147134
rect 505794 111454 506414 146898
rect 505794 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 506414 111454
rect 505794 111134 506414 111218
rect 505794 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 506414 111134
rect 505794 75454 506414 110898
rect 505794 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 506414 75454
rect 505794 75134 506414 75218
rect 505794 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 506414 75134
rect 505794 39454 506414 74898
rect 505794 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 506414 39454
rect 505794 39134 506414 39218
rect 505794 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 506414 39134
rect 505794 3454 506414 38898
rect 505794 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 506414 3454
rect 505794 3134 506414 3218
rect 505794 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 506414 3134
rect 505794 -346 506414 2898
rect 505794 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 506414 -346
rect 505794 -666 506414 -582
rect 505794 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 506414 -666
rect 505794 -1894 506414 -902
rect 509514 691174 510134 706202
rect 509514 690938 509546 691174
rect 509782 690938 509866 691174
rect 510102 690938 510134 691174
rect 509514 690854 510134 690938
rect 509514 690618 509546 690854
rect 509782 690618 509866 690854
rect 510102 690618 510134 690854
rect 509514 655174 510134 690618
rect 509514 654938 509546 655174
rect 509782 654938 509866 655174
rect 510102 654938 510134 655174
rect 509514 654854 510134 654938
rect 509514 654618 509546 654854
rect 509782 654618 509866 654854
rect 510102 654618 510134 654854
rect 509514 619174 510134 654618
rect 509514 618938 509546 619174
rect 509782 618938 509866 619174
rect 510102 618938 510134 619174
rect 509514 618854 510134 618938
rect 509514 618618 509546 618854
rect 509782 618618 509866 618854
rect 510102 618618 510134 618854
rect 509514 583174 510134 618618
rect 509514 582938 509546 583174
rect 509782 582938 509866 583174
rect 510102 582938 510134 583174
rect 509514 582854 510134 582938
rect 509514 582618 509546 582854
rect 509782 582618 509866 582854
rect 510102 582618 510134 582854
rect 509514 547174 510134 582618
rect 509514 546938 509546 547174
rect 509782 546938 509866 547174
rect 510102 546938 510134 547174
rect 509514 546854 510134 546938
rect 509514 546618 509546 546854
rect 509782 546618 509866 546854
rect 510102 546618 510134 546854
rect 509514 511174 510134 546618
rect 509514 510938 509546 511174
rect 509782 510938 509866 511174
rect 510102 510938 510134 511174
rect 509514 510854 510134 510938
rect 509514 510618 509546 510854
rect 509782 510618 509866 510854
rect 510102 510618 510134 510854
rect 509514 475174 510134 510618
rect 509514 474938 509546 475174
rect 509782 474938 509866 475174
rect 510102 474938 510134 475174
rect 509514 474854 510134 474938
rect 509514 474618 509546 474854
rect 509782 474618 509866 474854
rect 510102 474618 510134 474854
rect 509514 439174 510134 474618
rect 509514 438938 509546 439174
rect 509782 438938 509866 439174
rect 510102 438938 510134 439174
rect 509514 438854 510134 438938
rect 509514 438618 509546 438854
rect 509782 438618 509866 438854
rect 510102 438618 510134 438854
rect 509514 403174 510134 438618
rect 509514 402938 509546 403174
rect 509782 402938 509866 403174
rect 510102 402938 510134 403174
rect 509514 402854 510134 402938
rect 509514 402618 509546 402854
rect 509782 402618 509866 402854
rect 510102 402618 510134 402854
rect 509514 367174 510134 402618
rect 509514 366938 509546 367174
rect 509782 366938 509866 367174
rect 510102 366938 510134 367174
rect 509514 366854 510134 366938
rect 509514 366618 509546 366854
rect 509782 366618 509866 366854
rect 510102 366618 510134 366854
rect 509514 331174 510134 366618
rect 509514 330938 509546 331174
rect 509782 330938 509866 331174
rect 510102 330938 510134 331174
rect 509514 330854 510134 330938
rect 509514 330618 509546 330854
rect 509782 330618 509866 330854
rect 510102 330618 510134 330854
rect 509514 295174 510134 330618
rect 509514 294938 509546 295174
rect 509782 294938 509866 295174
rect 510102 294938 510134 295174
rect 509514 294854 510134 294938
rect 509514 294618 509546 294854
rect 509782 294618 509866 294854
rect 510102 294618 510134 294854
rect 509514 259174 510134 294618
rect 509514 258938 509546 259174
rect 509782 258938 509866 259174
rect 510102 258938 510134 259174
rect 509514 258854 510134 258938
rect 509514 258618 509546 258854
rect 509782 258618 509866 258854
rect 510102 258618 510134 258854
rect 509514 223174 510134 258618
rect 509514 222938 509546 223174
rect 509782 222938 509866 223174
rect 510102 222938 510134 223174
rect 509514 222854 510134 222938
rect 509514 222618 509546 222854
rect 509782 222618 509866 222854
rect 510102 222618 510134 222854
rect 509514 187174 510134 222618
rect 509514 186938 509546 187174
rect 509782 186938 509866 187174
rect 510102 186938 510134 187174
rect 509514 186854 510134 186938
rect 509514 186618 509546 186854
rect 509782 186618 509866 186854
rect 510102 186618 510134 186854
rect 509514 151174 510134 186618
rect 509514 150938 509546 151174
rect 509782 150938 509866 151174
rect 510102 150938 510134 151174
rect 509514 150854 510134 150938
rect 509514 150618 509546 150854
rect 509782 150618 509866 150854
rect 510102 150618 510134 150854
rect 509514 115174 510134 150618
rect 509514 114938 509546 115174
rect 509782 114938 509866 115174
rect 510102 114938 510134 115174
rect 509514 114854 510134 114938
rect 509514 114618 509546 114854
rect 509782 114618 509866 114854
rect 510102 114618 510134 114854
rect 509514 79174 510134 114618
rect 509514 78938 509546 79174
rect 509782 78938 509866 79174
rect 510102 78938 510134 79174
rect 509514 78854 510134 78938
rect 509514 78618 509546 78854
rect 509782 78618 509866 78854
rect 510102 78618 510134 78854
rect 509514 43174 510134 78618
rect 509514 42938 509546 43174
rect 509782 42938 509866 43174
rect 510102 42938 510134 43174
rect 509514 42854 510134 42938
rect 509514 42618 509546 42854
rect 509782 42618 509866 42854
rect 510102 42618 510134 42854
rect 509514 7174 510134 42618
rect 509514 6938 509546 7174
rect 509782 6938 509866 7174
rect 510102 6938 510134 7174
rect 509514 6854 510134 6938
rect 509514 6618 509546 6854
rect 509782 6618 509866 6854
rect 510102 6618 510134 6854
rect 509514 -2266 510134 6618
rect 509514 -2502 509546 -2266
rect 509782 -2502 509866 -2266
rect 510102 -2502 510134 -2266
rect 509514 -2586 510134 -2502
rect 509514 -2822 509546 -2586
rect 509782 -2822 509866 -2586
rect 510102 -2822 510134 -2586
rect 509514 -3814 510134 -2822
rect 513234 694894 513854 708122
rect 513234 694658 513266 694894
rect 513502 694658 513586 694894
rect 513822 694658 513854 694894
rect 513234 694574 513854 694658
rect 513234 694338 513266 694574
rect 513502 694338 513586 694574
rect 513822 694338 513854 694574
rect 513234 658894 513854 694338
rect 513234 658658 513266 658894
rect 513502 658658 513586 658894
rect 513822 658658 513854 658894
rect 513234 658574 513854 658658
rect 513234 658338 513266 658574
rect 513502 658338 513586 658574
rect 513822 658338 513854 658574
rect 513234 622894 513854 658338
rect 513234 622658 513266 622894
rect 513502 622658 513586 622894
rect 513822 622658 513854 622894
rect 513234 622574 513854 622658
rect 513234 622338 513266 622574
rect 513502 622338 513586 622574
rect 513822 622338 513854 622574
rect 513234 586894 513854 622338
rect 513234 586658 513266 586894
rect 513502 586658 513586 586894
rect 513822 586658 513854 586894
rect 513234 586574 513854 586658
rect 513234 586338 513266 586574
rect 513502 586338 513586 586574
rect 513822 586338 513854 586574
rect 513234 550894 513854 586338
rect 513234 550658 513266 550894
rect 513502 550658 513586 550894
rect 513822 550658 513854 550894
rect 513234 550574 513854 550658
rect 513234 550338 513266 550574
rect 513502 550338 513586 550574
rect 513822 550338 513854 550574
rect 513234 514894 513854 550338
rect 513234 514658 513266 514894
rect 513502 514658 513586 514894
rect 513822 514658 513854 514894
rect 513234 514574 513854 514658
rect 513234 514338 513266 514574
rect 513502 514338 513586 514574
rect 513822 514338 513854 514574
rect 513234 478894 513854 514338
rect 513234 478658 513266 478894
rect 513502 478658 513586 478894
rect 513822 478658 513854 478894
rect 513234 478574 513854 478658
rect 513234 478338 513266 478574
rect 513502 478338 513586 478574
rect 513822 478338 513854 478574
rect 513234 442894 513854 478338
rect 513234 442658 513266 442894
rect 513502 442658 513586 442894
rect 513822 442658 513854 442894
rect 513234 442574 513854 442658
rect 513234 442338 513266 442574
rect 513502 442338 513586 442574
rect 513822 442338 513854 442574
rect 513234 406894 513854 442338
rect 513234 406658 513266 406894
rect 513502 406658 513586 406894
rect 513822 406658 513854 406894
rect 513234 406574 513854 406658
rect 513234 406338 513266 406574
rect 513502 406338 513586 406574
rect 513822 406338 513854 406574
rect 513234 370894 513854 406338
rect 513234 370658 513266 370894
rect 513502 370658 513586 370894
rect 513822 370658 513854 370894
rect 513234 370574 513854 370658
rect 513234 370338 513266 370574
rect 513502 370338 513586 370574
rect 513822 370338 513854 370574
rect 513234 334894 513854 370338
rect 513234 334658 513266 334894
rect 513502 334658 513586 334894
rect 513822 334658 513854 334894
rect 513234 334574 513854 334658
rect 513234 334338 513266 334574
rect 513502 334338 513586 334574
rect 513822 334338 513854 334574
rect 513234 298894 513854 334338
rect 513234 298658 513266 298894
rect 513502 298658 513586 298894
rect 513822 298658 513854 298894
rect 513234 298574 513854 298658
rect 513234 298338 513266 298574
rect 513502 298338 513586 298574
rect 513822 298338 513854 298574
rect 513234 262894 513854 298338
rect 513234 262658 513266 262894
rect 513502 262658 513586 262894
rect 513822 262658 513854 262894
rect 513234 262574 513854 262658
rect 513234 262338 513266 262574
rect 513502 262338 513586 262574
rect 513822 262338 513854 262574
rect 513234 226894 513854 262338
rect 513234 226658 513266 226894
rect 513502 226658 513586 226894
rect 513822 226658 513854 226894
rect 513234 226574 513854 226658
rect 513234 226338 513266 226574
rect 513502 226338 513586 226574
rect 513822 226338 513854 226574
rect 513234 190894 513854 226338
rect 513234 190658 513266 190894
rect 513502 190658 513586 190894
rect 513822 190658 513854 190894
rect 513234 190574 513854 190658
rect 513234 190338 513266 190574
rect 513502 190338 513586 190574
rect 513822 190338 513854 190574
rect 513234 154894 513854 190338
rect 513234 154658 513266 154894
rect 513502 154658 513586 154894
rect 513822 154658 513854 154894
rect 513234 154574 513854 154658
rect 513234 154338 513266 154574
rect 513502 154338 513586 154574
rect 513822 154338 513854 154574
rect 513234 118894 513854 154338
rect 513234 118658 513266 118894
rect 513502 118658 513586 118894
rect 513822 118658 513854 118894
rect 513234 118574 513854 118658
rect 513234 118338 513266 118574
rect 513502 118338 513586 118574
rect 513822 118338 513854 118574
rect 513234 82894 513854 118338
rect 513234 82658 513266 82894
rect 513502 82658 513586 82894
rect 513822 82658 513854 82894
rect 513234 82574 513854 82658
rect 513234 82338 513266 82574
rect 513502 82338 513586 82574
rect 513822 82338 513854 82574
rect 513234 46894 513854 82338
rect 513234 46658 513266 46894
rect 513502 46658 513586 46894
rect 513822 46658 513854 46894
rect 513234 46574 513854 46658
rect 513234 46338 513266 46574
rect 513502 46338 513586 46574
rect 513822 46338 513854 46574
rect 513234 10894 513854 46338
rect 513234 10658 513266 10894
rect 513502 10658 513586 10894
rect 513822 10658 513854 10894
rect 513234 10574 513854 10658
rect 513234 10338 513266 10574
rect 513502 10338 513586 10574
rect 513822 10338 513854 10574
rect 513234 -4186 513854 10338
rect 513234 -4422 513266 -4186
rect 513502 -4422 513586 -4186
rect 513822 -4422 513854 -4186
rect 513234 -4506 513854 -4422
rect 513234 -4742 513266 -4506
rect 513502 -4742 513586 -4506
rect 513822 -4742 513854 -4506
rect 513234 -5734 513854 -4742
rect 516954 698614 517574 710042
rect 534954 711558 535574 711590
rect 534954 711322 534986 711558
rect 535222 711322 535306 711558
rect 535542 711322 535574 711558
rect 534954 711238 535574 711322
rect 534954 711002 534986 711238
rect 535222 711002 535306 711238
rect 535542 711002 535574 711238
rect 531234 709638 531854 709670
rect 531234 709402 531266 709638
rect 531502 709402 531586 709638
rect 531822 709402 531854 709638
rect 531234 709318 531854 709402
rect 531234 709082 531266 709318
rect 531502 709082 531586 709318
rect 531822 709082 531854 709318
rect 527514 707718 528134 707750
rect 527514 707482 527546 707718
rect 527782 707482 527866 707718
rect 528102 707482 528134 707718
rect 527514 707398 528134 707482
rect 527514 707162 527546 707398
rect 527782 707162 527866 707398
rect 528102 707162 528134 707398
rect 516954 698378 516986 698614
rect 517222 698378 517306 698614
rect 517542 698378 517574 698614
rect 516954 698294 517574 698378
rect 516954 698058 516986 698294
rect 517222 698058 517306 698294
rect 517542 698058 517574 698294
rect 516954 662614 517574 698058
rect 516954 662378 516986 662614
rect 517222 662378 517306 662614
rect 517542 662378 517574 662614
rect 516954 662294 517574 662378
rect 516954 662058 516986 662294
rect 517222 662058 517306 662294
rect 517542 662058 517574 662294
rect 516954 626614 517574 662058
rect 516954 626378 516986 626614
rect 517222 626378 517306 626614
rect 517542 626378 517574 626614
rect 516954 626294 517574 626378
rect 516954 626058 516986 626294
rect 517222 626058 517306 626294
rect 517542 626058 517574 626294
rect 516954 590614 517574 626058
rect 516954 590378 516986 590614
rect 517222 590378 517306 590614
rect 517542 590378 517574 590614
rect 516954 590294 517574 590378
rect 516954 590058 516986 590294
rect 517222 590058 517306 590294
rect 517542 590058 517574 590294
rect 516954 554614 517574 590058
rect 516954 554378 516986 554614
rect 517222 554378 517306 554614
rect 517542 554378 517574 554614
rect 516954 554294 517574 554378
rect 516954 554058 516986 554294
rect 517222 554058 517306 554294
rect 517542 554058 517574 554294
rect 516954 518614 517574 554058
rect 516954 518378 516986 518614
rect 517222 518378 517306 518614
rect 517542 518378 517574 518614
rect 516954 518294 517574 518378
rect 516954 518058 516986 518294
rect 517222 518058 517306 518294
rect 517542 518058 517574 518294
rect 516954 482614 517574 518058
rect 516954 482378 516986 482614
rect 517222 482378 517306 482614
rect 517542 482378 517574 482614
rect 516954 482294 517574 482378
rect 516954 482058 516986 482294
rect 517222 482058 517306 482294
rect 517542 482058 517574 482294
rect 516954 446614 517574 482058
rect 516954 446378 516986 446614
rect 517222 446378 517306 446614
rect 517542 446378 517574 446614
rect 516954 446294 517574 446378
rect 516954 446058 516986 446294
rect 517222 446058 517306 446294
rect 517542 446058 517574 446294
rect 516954 410614 517574 446058
rect 516954 410378 516986 410614
rect 517222 410378 517306 410614
rect 517542 410378 517574 410614
rect 516954 410294 517574 410378
rect 516954 410058 516986 410294
rect 517222 410058 517306 410294
rect 517542 410058 517574 410294
rect 516954 374614 517574 410058
rect 516954 374378 516986 374614
rect 517222 374378 517306 374614
rect 517542 374378 517574 374614
rect 516954 374294 517574 374378
rect 516954 374058 516986 374294
rect 517222 374058 517306 374294
rect 517542 374058 517574 374294
rect 516954 338614 517574 374058
rect 516954 338378 516986 338614
rect 517222 338378 517306 338614
rect 517542 338378 517574 338614
rect 516954 338294 517574 338378
rect 516954 338058 516986 338294
rect 517222 338058 517306 338294
rect 517542 338058 517574 338294
rect 516954 302614 517574 338058
rect 516954 302378 516986 302614
rect 517222 302378 517306 302614
rect 517542 302378 517574 302614
rect 516954 302294 517574 302378
rect 516954 302058 516986 302294
rect 517222 302058 517306 302294
rect 517542 302058 517574 302294
rect 516954 266614 517574 302058
rect 516954 266378 516986 266614
rect 517222 266378 517306 266614
rect 517542 266378 517574 266614
rect 516954 266294 517574 266378
rect 516954 266058 516986 266294
rect 517222 266058 517306 266294
rect 517542 266058 517574 266294
rect 516954 230614 517574 266058
rect 516954 230378 516986 230614
rect 517222 230378 517306 230614
rect 517542 230378 517574 230614
rect 516954 230294 517574 230378
rect 516954 230058 516986 230294
rect 517222 230058 517306 230294
rect 517542 230058 517574 230294
rect 516954 194614 517574 230058
rect 516954 194378 516986 194614
rect 517222 194378 517306 194614
rect 517542 194378 517574 194614
rect 516954 194294 517574 194378
rect 516954 194058 516986 194294
rect 517222 194058 517306 194294
rect 517542 194058 517574 194294
rect 516954 158614 517574 194058
rect 516954 158378 516986 158614
rect 517222 158378 517306 158614
rect 517542 158378 517574 158614
rect 516954 158294 517574 158378
rect 516954 158058 516986 158294
rect 517222 158058 517306 158294
rect 517542 158058 517574 158294
rect 516954 122614 517574 158058
rect 516954 122378 516986 122614
rect 517222 122378 517306 122614
rect 517542 122378 517574 122614
rect 516954 122294 517574 122378
rect 516954 122058 516986 122294
rect 517222 122058 517306 122294
rect 517542 122058 517574 122294
rect 516954 86614 517574 122058
rect 516954 86378 516986 86614
rect 517222 86378 517306 86614
rect 517542 86378 517574 86614
rect 516954 86294 517574 86378
rect 516954 86058 516986 86294
rect 517222 86058 517306 86294
rect 517542 86058 517574 86294
rect 516954 50614 517574 86058
rect 516954 50378 516986 50614
rect 517222 50378 517306 50614
rect 517542 50378 517574 50614
rect 516954 50294 517574 50378
rect 516954 50058 516986 50294
rect 517222 50058 517306 50294
rect 517542 50058 517574 50294
rect 516954 14614 517574 50058
rect 516954 14378 516986 14614
rect 517222 14378 517306 14614
rect 517542 14378 517574 14614
rect 516954 14294 517574 14378
rect 516954 14058 516986 14294
rect 517222 14058 517306 14294
rect 517542 14058 517574 14294
rect 498954 -7302 498986 -7066
rect 499222 -7302 499306 -7066
rect 499542 -7302 499574 -7066
rect 498954 -7386 499574 -7302
rect 498954 -7622 498986 -7386
rect 499222 -7622 499306 -7386
rect 499542 -7622 499574 -7386
rect 498954 -7654 499574 -7622
rect 516954 -6106 517574 14058
rect 523794 705798 524414 705830
rect 523794 705562 523826 705798
rect 524062 705562 524146 705798
rect 524382 705562 524414 705798
rect 523794 705478 524414 705562
rect 523794 705242 523826 705478
rect 524062 705242 524146 705478
rect 524382 705242 524414 705478
rect 523794 669454 524414 705242
rect 523794 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 524414 669454
rect 523794 669134 524414 669218
rect 523794 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 524414 669134
rect 523794 633454 524414 668898
rect 523794 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 524414 633454
rect 523794 633134 524414 633218
rect 523794 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 524414 633134
rect 523794 597454 524414 632898
rect 523794 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 524414 597454
rect 523794 597134 524414 597218
rect 523794 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 524414 597134
rect 523794 561454 524414 596898
rect 523794 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 524414 561454
rect 523794 561134 524414 561218
rect 523794 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 524414 561134
rect 523794 525454 524414 560898
rect 523794 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 524414 525454
rect 523794 525134 524414 525218
rect 523794 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 524414 525134
rect 523794 489454 524414 524898
rect 523794 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 524414 489454
rect 523794 489134 524414 489218
rect 523794 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 524414 489134
rect 523794 453454 524414 488898
rect 523794 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 524414 453454
rect 523794 453134 524414 453218
rect 523794 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 524414 453134
rect 523794 417454 524414 452898
rect 523794 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 524414 417454
rect 523794 417134 524414 417218
rect 523794 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 524414 417134
rect 523794 381454 524414 416898
rect 523794 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 524414 381454
rect 523794 381134 524414 381218
rect 523794 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 524414 381134
rect 523794 345454 524414 380898
rect 523794 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 524414 345454
rect 523794 345134 524414 345218
rect 523794 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 524414 345134
rect 523794 309454 524414 344898
rect 523794 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 524414 309454
rect 523794 309134 524414 309218
rect 523794 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 524414 309134
rect 523794 273454 524414 308898
rect 523794 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 524414 273454
rect 523794 273134 524414 273218
rect 523794 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 524414 273134
rect 523794 237454 524414 272898
rect 523794 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 524414 237454
rect 523794 237134 524414 237218
rect 523794 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 524414 237134
rect 523794 201454 524414 236898
rect 523794 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 524414 201454
rect 523794 201134 524414 201218
rect 523794 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 524414 201134
rect 523794 165454 524414 200898
rect 523794 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 524414 165454
rect 523794 165134 524414 165218
rect 523794 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 524414 165134
rect 523794 129454 524414 164898
rect 523794 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 524414 129454
rect 523794 129134 524414 129218
rect 523794 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 524414 129134
rect 523794 93454 524414 128898
rect 523794 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 524414 93454
rect 523794 93134 524414 93218
rect 523794 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 524414 93134
rect 523794 57454 524414 92898
rect 523794 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 524414 57454
rect 523794 57134 524414 57218
rect 523794 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 524414 57134
rect 523794 21454 524414 56898
rect 523794 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 524414 21454
rect 523794 21134 524414 21218
rect 523794 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 524414 21134
rect 523794 -1306 524414 20898
rect 523794 -1542 523826 -1306
rect 524062 -1542 524146 -1306
rect 524382 -1542 524414 -1306
rect 523794 -1626 524414 -1542
rect 523794 -1862 523826 -1626
rect 524062 -1862 524146 -1626
rect 524382 -1862 524414 -1626
rect 523794 -1894 524414 -1862
rect 527514 673174 528134 707162
rect 527514 672938 527546 673174
rect 527782 672938 527866 673174
rect 528102 672938 528134 673174
rect 527514 672854 528134 672938
rect 527514 672618 527546 672854
rect 527782 672618 527866 672854
rect 528102 672618 528134 672854
rect 527514 637174 528134 672618
rect 527514 636938 527546 637174
rect 527782 636938 527866 637174
rect 528102 636938 528134 637174
rect 527514 636854 528134 636938
rect 527514 636618 527546 636854
rect 527782 636618 527866 636854
rect 528102 636618 528134 636854
rect 527514 601174 528134 636618
rect 527514 600938 527546 601174
rect 527782 600938 527866 601174
rect 528102 600938 528134 601174
rect 527514 600854 528134 600938
rect 527514 600618 527546 600854
rect 527782 600618 527866 600854
rect 528102 600618 528134 600854
rect 527514 565174 528134 600618
rect 527514 564938 527546 565174
rect 527782 564938 527866 565174
rect 528102 564938 528134 565174
rect 527514 564854 528134 564938
rect 527514 564618 527546 564854
rect 527782 564618 527866 564854
rect 528102 564618 528134 564854
rect 527514 529174 528134 564618
rect 527514 528938 527546 529174
rect 527782 528938 527866 529174
rect 528102 528938 528134 529174
rect 527514 528854 528134 528938
rect 527514 528618 527546 528854
rect 527782 528618 527866 528854
rect 528102 528618 528134 528854
rect 527514 493174 528134 528618
rect 527514 492938 527546 493174
rect 527782 492938 527866 493174
rect 528102 492938 528134 493174
rect 527514 492854 528134 492938
rect 527514 492618 527546 492854
rect 527782 492618 527866 492854
rect 528102 492618 528134 492854
rect 527514 457174 528134 492618
rect 527514 456938 527546 457174
rect 527782 456938 527866 457174
rect 528102 456938 528134 457174
rect 527514 456854 528134 456938
rect 527514 456618 527546 456854
rect 527782 456618 527866 456854
rect 528102 456618 528134 456854
rect 527514 421174 528134 456618
rect 527514 420938 527546 421174
rect 527782 420938 527866 421174
rect 528102 420938 528134 421174
rect 527514 420854 528134 420938
rect 527514 420618 527546 420854
rect 527782 420618 527866 420854
rect 528102 420618 528134 420854
rect 527514 385174 528134 420618
rect 527514 384938 527546 385174
rect 527782 384938 527866 385174
rect 528102 384938 528134 385174
rect 527514 384854 528134 384938
rect 527514 384618 527546 384854
rect 527782 384618 527866 384854
rect 528102 384618 528134 384854
rect 527514 349174 528134 384618
rect 527514 348938 527546 349174
rect 527782 348938 527866 349174
rect 528102 348938 528134 349174
rect 527514 348854 528134 348938
rect 527514 348618 527546 348854
rect 527782 348618 527866 348854
rect 528102 348618 528134 348854
rect 527514 313174 528134 348618
rect 527514 312938 527546 313174
rect 527782 312938 527866 313174
rect 528102 312938 528134 313174
rect 527514 312854 528134 312938
rect 527514 312618 527546 312854
rect 527782 312618 527866 312854
rect 528102 312618 528134 312854
rect 527514 277174 528134 312618
rect 527514 276938 527546 277174
rect 527782 276938 527866 277174
rect 528102 276938 528134 277174
rect 527514 276854 528134 276938
rect 527514 276618 527546 276854
rect 527782 276618 527866 276854
rect 528102 276618 528134 276854
rect 527514 241174 528134 276618
rect 527514 240938 527546 241174
rect 527782 240938 527866 241174
rect 528102 240938 528134 241174
rect 527514 240854 528134 240938
rect 527514 240618 527546 240854
rect 527782 240618 527866 240854
rect 528102 240618 528134 240854
rect 527514 205174 528134 240618
rect 527514 204938 527546 205174
rect 527782 204938 527866 205174
rect 528102 204938 528134 205174
rect 527514 204854 528134 204938
rect 527514 204618 527546 204854
rect 527782 204618 527866 204854
rect 528102 204618 528134 204854
rect 527514 169174 528134 204618
rect 527514 168938 527546 169174
rect 527782 168938 527866 169174
rect 528102 168938 528134 169174
rect 527514 168854 528134 168938
rect 527514 168618 527546 168854
rect 527782 168618 527866 168854
rect 528102 168618 528134 168854
rect 527514 133174 528134 168618
rect 527514 132938 527546 133174
rect 527782 132938 527866 133174
rect 528102 132938 528134 133174
rect 527514 132854 528134 132938
rect 527514 132618 527546 132854
rect 527782 132618 527866 132854
rect 528102 132618 528134 132854
rect 527514 97174 528134 132618
rect 527514 96938 527546 97174
rect 527782 96938 527866 97174
rect 528102 96938 528134 97174
rect 527514 96854 528134 96938
rect 527514 96618 527546 96854
rect 527782 96618 527866 96854
rect 528102 96618 528134 96854
rect 527514 61174 528134 96618
rect 527514 60938 527546 61174
rect 527782 60938 527866 61174
rect 528102 60938 528134 61174
rect 527514 60854 528134 60938
rect 527514 60618 527546 60854
rect 527782 60618 527866 60854
rect 528102 60618 528134 60854
rect 527514 25174 528134 60618
rect 527514 24938 527546 25174
rect 527782 24938 527866 25174
rect 528102 24938 528134 25174
rect 527514 24854 528134 24938
rect 527514 24618 527546 24854
rect 527782 24618 527866 24854
rect 528102 24618 528134 24854
rect 527514 -3226 528134 24618
rect 527514 -3462 527546 -3226
rect 527782 -3462 527866 -3226
rect 528102 -3462 528134 -3226
rect 527514 -3546 528134 -3462
rect 527514 -3782 527546 -3546
rect 527782 -3782 527866 -3546
rect 528102 -3782 528134 -3546
rect 527514 -3814 528134 -3782
rect 531234 676894 531854 709082
rect 531234 676658 531266 676894
rect 531502 676658 531586 676894
rect 531822 676658 531854 676894
rect 531234 676574 531854 676658
rect 531234 676338 531266 676574
rect 531502 676338 531586 676574
rect 531822 676338 531854 676574
rect 531234 640894 531854 676338
rect 531234 640658 531266 640894
rect 531502 640658 531586 640894
rect 531822 640658 531854 640894
rect 531234 640574 531854 640658
rect 531234 640338 531266 640574
rect 531502 640338 531586 640574
rect 531822 640338 531854 640574
rect 531234 604894 531854 640338
rect 531234 604658 531266 604894
rect 531502 604658 531586 604894
rect 531822 604658 531854 604894
rect 531234 604574 531854 604658
rect 531234 604338 531266 604574
rect 531502 604338 531586 604574
rect 531822 604338 531854 604574
rect 531234 568894 531854 604338
rect 531234 568658 531266 568894
rect 531502 568658 531586 568894
rect 531822 568658 531854 568894
rect 531234 568574 531854 568658
rect 531234 568338 531266 568574
rect 531502 568338 531586 568574
rect 531822 568338 531854 568574
rect 531234 532894 531854 568338
rect 531234 532658 531266 532894
rect 531502 532658 531586 532894
rect 531822 532658 531854 532894
rect 531234 532574 531854 532658
rect 531234 532338 531266 532574
rect 531502 532338 531586 532574
rect 531822 532338 531854 532574
rect 531234 496894 531854 532338
rect 531234 496658 531266 496894
rect 531502 496658 531586 496894
rect 531822 496658 531854 496894
rect 531234 496574 531854 496658
rect 531234 496338 531266 496574
rect 531502 496338 531586 496574
rect 531822 496338 531854 496574
rect 531234 460894 531854 496338
rect 531234 460658 531266 460894
rect 531502 460658 531586 460894
rect 531822 460658 531854 460894
rect 531234 460574 531854 460658
rect 531234 460338 531266 460574
rect 531502 460338 531586 460574
rect 531822 460338 531854 460574
rect 531234 424894 531854 460338
rect 531234 424658 531266 424894
rect 531502 424658 531586 424894
rect 531822 424658 531854 424894
rect 531234 424574 531854 424658
rect 531234 424338 531266 424574
rect 531502 424338 531586 424574
rect 531822 424338 531854 424574
rect 531234 388894 531854 424338
rect 531234 388658 531266 388894
rect 531502 388658 531586 388894
rect 531822 388658 531854 388894
rect 531234 388574 531854 388658
rect 531234 388338 531266 388574
rect 531502 388338 531586 388574
rect 531822 388338 531854 388574
rect 531234 352894 531854 388338
rect 531234 352658 531266 352894
rect 531502 352658 531586 352894
rect 531822 352658 531854 352894
rect 531234 352574 531854 352658
rect 531234 352338 531266 352574
rect 531502 352338 531586 352574
rect 531822 352338 531854 352574
rect 531234 316894 531854 352338
rect 531234 316658 531266 316894
rect 531502 316658 531586 316894
rect 531822 316658 531854 316894
rect 531234 316574 531854 316658
rect 531234 316338 531266 316574
rect 531502 316338 531586 316574
rect 531822 316338 531854 316574
rect 531234 280894 531854 316338
rect 531234 280658 531266 280894
rect 531502 280658 531586 280894
rect 531822 280658 531854 280894
rect 531234 280574 531854 280658
rect 531234 280338 531266 280574
rect 531502 280338 531586 280574
rect 531822 280338 531854 280574
rect 531234 244894 531854 280338
rect 531234 244658 531266 244894
rect 531502 244658 531586 244894
rect 531822 244658 531854 244894
rect 531234 244574 531854 244658
rect 531234 244338 531266 244574
rect 531502 244338 531586 244574
rect 531822 244338 531854 244574
rect 531234 208894 531854 244338
rect 531234 208658 531266 208894
rect 531502 208658 531586 208894
rect 531822 208658 531854 208894
rect 531234 208574 531854 208658
rect 531234 208338 531266 208574
rect 531502 208338 531586 208574
rect 531822 208338 531854 208574
rect 531234 172894 531854 208338
rect 531234 172658 531266 172894
rect 531502 172658 531586 172894
rect 531822 172658 531854 172894
rect 531234 172574 531854 172658
rect 531234 172338 531266 172574
rect 531502 172338 531586 172574
rect 531822 172338 531854 172574
rect 531234 136894 531854 172338
rect 531234 136658 531266 136894
rect 531502 136658 531586 136894
rect 531822 136658 531854 136894
rect 531234 136574 531854 136658
rect 531234 136338 531266 136574
rect 531502 136338 531586 136574
rect 531822 136338 531854 136574
rect 531234 100894 531854 136338
rect 531234 100658 531266 100894
rect 531502 100658 531586 100894
rect 531822 100658 531854 100894
rect 531234 100574 531854 100658
rect 531234 100338 531266 100574
rect 531502 100338 531586 100574
rect 531822 100338 531854 100574
rect 531234 64894 531854 100338
rect 531234 64658 531266 64894
rect 531502 64658 531586 64894
rect 531822 64658 531854 64894
rect 531234 64574 531854 64658
rect 531234 64338 531266 64574
rect 531502 64338 531586 64574
rect 531822 64338 531854 64574
rect 531234 28894 531854 64338
rect 531234 28658 531266 28894
rect 531502 28658 531586 28894
rect 531822 28658 531854 28894
rect 531234 28574 531854 28658
rect 531234 28338 531266 28574
rect 531502 28338 531586 28574
rect 531822 28338 531854 28574
rect 531234 -5146 531854 28338
rect 531234 -5382 531266 -5146
rect 531502 -5382 531586 -5146
rect 531822 -5382 531854 -5146
rect 531234 -5466 531854 -5382
rect 531234 -5702 531266 -5466
rect 531502 -5702 531586 -5466
rect 531822 -5702 531854 -5466
rect 531234 -5734 531854 -5702
rect 534954 680614 535574 711002
rect 552954 710598 553574 711590
rect 552954 710362 552986 710598
rect 553222 710362 553306 710598
rect 553542 710362 553574 710598
rect 552954 710278 553574 710362
rect 552954 710042 552986 710278
rect 553222 710042 553306 710278
rect 553542 710042 553574 710278
rect 549234 708678 549854 709670
rect 549234 708442 549266 708678
rect 549502 708442 549586 708678
rect 549822 708442 549854 708678
rect 549234 708358 549854 708442
rect 549234 708122 549266 708358
rect 549502 708122 549586 708358
rect 549822 708122 549854 708358
rect 545514 706758 546134 707750
rect 545514 706522 545546 706758
rect 545782 706522 545866 706758
rect 546102 706522 546134 706758
rect 545514 706438 546134 706522
rect 545514 706202 545546 706438
rect 545782 706202 545866 706438
rect 546102 706202 546134 706438
rect 534954 680378 534986 680614
rect 535222 680378 535306 680614
rect 535542 680378 535574 680614
rect 534954 680294 535574 680378
rect 534954 680058 534986 680294
rect 535222 680058 535306 680294
rect 535542 680058 535574 680294
rect 534954 644614 535574 680058
rect 534954 644378 534986 644614
rect 535222 644378 535306 644614
rect 535542 644378 535574 644614
rect 534954 644294 535574 644378
rect 534954 644058 534986 644294
rect 535222 644058 535306 644294
rect 535542 644058 535574 644294
rect 534954 608614 535574 644058
rect 534954 608378 534986 608614
rect 535222 608378 535306 608614
rect 535542 608378 535574 608614
rect 534954 608294 535574 608378
rect 534954 608058 534986 608294
rect 535222 608058 535306 608294
rect 535542 608058 535574 608294
rect 534954 572614 535574 608058
rect 534954 572378 534986 572614
rect 535222 572378 535306 572614
rect 535542 572378 535574 572614
rect 534954 572294 535574 572378
rect 534954 572058 534986 572294
rect 535222 572058 535306 572294
rect 535542 572058 535574 572294
rect 534954 536614 535574 572058
rect 534954 536378 534986 536614
rect 535222 536378 535306 536614
rect 535542 536378 535574 536614
rect 534954 536294 535574 536378
rect 534954 536058 534986 536294
rect 535222 536058 535306 536294
rect 535542 536058 535574 536294
rect 534954 500614 535574 536058
rect 534954 500378 534986 500614
rect 535222 500378 535306 500614
rect 535542 500378 535574 500614
rect 534954 500294 535574 500378
rect 534954 500058 534986 500294
rect 535222 500058 535306 500294
rect 535542 500058 535574 500294
rect 534954 464614 535574 500058
rect 534954 464378 534986 464614
rect 535222 464378 535306 464614
rect 535542 464378 535574 464614
rect 534954 464294 535574 464378
rect 534954 464058 534986 464294
rect 535222 464058 535306 464294
rect 535542 464058 535574 464294
rect 534954 428614 535574 464058
rect 534954 428378 534986 428614
rect 535222 428378 535306 428614
rect 535542 428378 535574 428614
rect 534954 428294 535574 428378
rect 534954 428058 534986 428294
rect 535222 428058 535306 428294
rect 535542 428058 535574 428294
rect 534954 392614 535574 428058
rect 534954 392378 534986 392614
rect 535222 392378 535306 392614
rect 535542 392378 535574 392614
rect 534954 392294 535574 392378
rect 534954 392058 534986 392294
rect 535222 392058 535306 392294
rect 535542 392058 535574 392294
rect 534954 356614 535574 392058
rect 534954 356378 534986 356614
rect 535222 356378 535306 356614
rect 535542 356378 535574 356614
rect 534954 356294 535574 356378
rect 534954 356058 534986 356294
rect 535222 356058 535306 356294
rect 535542 356058 535574 356294
rect 534954 320614 535574 356058
rect 534954 320378 534986 320614
rect 535222 320378 535306 320614
rect 535542 320378 535574 320614
rect 534954 320294 535574 320378
rect 534954 320058 534986 320294
rect 535222 320058 535306 320294
rect 535542 320058 535574 320294
rect 534954 284614 535574 320058
rect 534954 284378 534986 284614
rect 535222 284378 535306 284614
rect 535542 284378 535574 284614
rect 534954 284294 535574 284378
rect 534954 284058 534986 284294
rect 535222 284058 535306 284294
rect 535542 284058 535574 284294
rect 534954 248614 535574 284058
rect 534954 248378 534986 248614
rect 535222 248378 535306 248614
rect 535542 248378 535574 248614
rect 534954 248294 535574 248378
rect 534954 248058 534986 248294
rect 535222 248058 535306 248294
rect 535542 248058 535574 248294
rect 534954 212614 535574 248058
rect 534954 212378 534986 212614
rect 535222 212378 535306 212614
rect 535542 212378 535574 212614
rect 534954 212294 535574 212378
rect 534954 212058 534986 212294
rect 535222 212058 535306 212294
rect 535542 212058 535574 212294
rect 534954 176614 535574 212058
rect 534954 176378 534986 176614
rect 535222 176378 535306 176614
rect 535542 176378 535574 176614
rect 534954 176294 535574 176378
rect 534954 176058 534986 176294
rect 535222 176058 535306 176294
rect 535542 176058 535574 176294
rect 534954 140614 535574 176058
rect 534954 140378 534986 140614
rect 535222 140378 535306 140614
rect 535542 140378 535574 140614
rect 534954 140294 535574 140378
rect 534954 140058 534986 140294
rect 535222 140058 535306 140294
rect 535542 140058 535574 140294
rect 534954 104614 535574 140058
rect 534954 104378 534986 104614
rect 535222 104378 535306 104614
rect 535542 104378 535574 104614
rect 534954 104294 535574 104378
rect 534954 104058 534986 104294
rect 535222 104058 535306 104294
rect 535542 104058 535574 104294
rect 534954 68614 535574 104058
rect 534954 68378 534986 68614
rect 535222 68378 535306 68614
rect 535542 68378 535574 68614
rect 534954 68294 535574 68378
rect 534954 68058 534986 68294
rect 535222 68058 535306 68294
rect 535542 68058 535574 68294
rect 534954 32614 535574 68058
rect 534954 32378 534986 32614
rect 535222 32378 535306 32614
rect 535542 32378 535574 32614
rect 534954 32294 535574 32378
rect 534954 32058 534986 32294
rect 535222 32058 535306 32294
rect 535542 32058 535574 32294
rect 516954 -6342 516986 -6106
rect 517222 -6342 517306 -6106
rect 517542 -6342 517574 -6106
rect 516954 -6426 517574 -6342
rect 516954 -6662 516986 -6426
rect 517222 -6662 517306 -6426
rect 517542 -6662 517574 -6426
rect 516954 -7654 517574 -6662
rect 534954 -7066 535574 32058
rect 541794 704838 542414 705830
rect 541794 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 542414 704838
rect 541794 704518 542414 704602
rect 541794 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 542414 704518
rect 541794 687454 542414 704282
rect 541794 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 542414 687454
rect 541794 687134 542414 687218
rect 541794 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 542414 687134
rect 541794 651454 542414 686898
rect 541794 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 542414 651454
rect 541794 651134 542414 651218
rect 541794 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 542414 651134
rect 541794 615454 542414 650898
rect 541794 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 542414 615454
rect 541794 615134 542414 615218
rect 541794 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 542414 615134
rect 541794 579454 542414 614898
rect 541794 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 542414 579454
rect 541794 579134 542414 579218
rect 541794 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 542414 579134
rect 541794 543454 542414 578898
rect 541794 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 542414 543454
rect 541794 543134 542414 543218
rect 541794 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 542414 543134
rect 541794 507454 542414 542898
rect 541794 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 542414 507454
rect 541794 507134 542414 507218
rect 541794 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 542414 507134
rect 541794 471454 542414 506898
rect 541794 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 542414 471454
rect 541794 471134 542414 471218
rect 541794 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 542414 471134
rect 541794 435454 542414 470898
rect 541794 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 542414 435454
rect 541794 435134 542414 435218
rect 541794 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 542414 435134
rect 541794 399454 542414 434898
rect 541794 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 542414 399454
rect 541794 399134 542414 399218
rect 541794 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 542414 399134
rect 541794 363454 542414 398898
rect 541794 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 542414 363454
rect 541794 363134 542414 363218
rect 541794 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 542414 363134
rect 541794 327454 542414 362898
rect 541794 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 542414 327454
rect 541794 327134 542414 327218
rect 541794 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 542414 327134
rect 541794 291454 542414 326898
rect 541794 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 542414 291454
rect 541794 291134 542414 291218
rect 541794 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 542414 291134
rect 541794 255454 542414 290898
rect 541794 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 542414 255454
rect 541794 255134 542414 255218
rect 541794 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 542414 255134
rect 541794 219454 542414 254898
rect 541794 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 542414 219454
rect 541794 219134 542414 219218
rect 541794 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 542414 219134
rect 541794 183454 542414 218898
rect 541794 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 542414 183454
rect 541794 183134 542414 183218
rect 541794 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 542414 183134
rect 541794 147454 542414 182898
rect 541794 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 542414 147454
rect 541794 147134 542414 147218
rect 541794 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 542414 147134
rect 541794 111454 542414 146898
rect 541794 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 542414 111454
rect 541794 111134 542414 111218
rect 541794 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 542414 111134
rect 541794 75454 542414 110898
rect 541794 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 542414 75454
rect 541794 75134 542414 75218
rect 541794 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 542414 75134
rect 541794 39454 542414 74898
rect 541794 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 542414 39454
rect 541794 39134 542414 39218
rect 541794 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 542414 39134
rect 541794 3454 542414 38898
rect 541794 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 542414 3454
rect 541794 3134 542414 3218
rect 541794 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 542414 3134
rect 541794 -346 542414 2898
rect 541794 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 542414 -346
rect 541794 -666 542414 -582
rect 541794 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 542414 -666
rect 541794 -1894 542414 -902
rect 545514 691174 546134 706202
rect 545514 690938 545546 691174
rect 545782 690938 545866 691174
rect 546102 690938 546134 691174
rect 545514 690854 546134 690938
rect 545514 690618 545546 690854
rect 545782 690618 545866 690854
rect 546102 690618 546134 690854
rect 545514 655174 546134 690618
rect 545514 654938 545546 655174
rect 545782 654938 545866 655174
rect 546102 654938 546134 655174
rect 545514 654854 546134 654938
rect 545514 654618 545546 654854
rect 545782 654618 545866 654854
rect 546102 654618 546134 654854
rect 545514 619174 546134 654618
rect 545514 618938 545546 619174
rect 545782 618938 545866 619174
rect 546102 618938 546134 619174
rect 545514 618854 546134 618938
rect 545514 618618 545546 618854
rect 545782 618618 545866 618854
rect 546102 618618 546134 618854
rect 545514 583174 546134 618618
rect 545514 582938 545546 583174
rect 545782 582938 545866 583174
rect 546102 582938 546134 583174
rect 545514 582854 546134 582938
rect 545514 582618 545546 582854
rect 545782 582618 545866 582854
rect 546102 582618 546134 582854
rect 545514 547174 546134 582618
rect 545514 546938 545546 547174
rect 545782 546938 545866 547174
rect 546102 546938 546134 547174
rect 545514 546854 546134 546938
rect 545514 546618 545546 546854
rect 545782 546618 545866 546854
rect 546102 546618 546134 546854
rect 545514 511174 546134 546618
rect 545514 510938 545546 511174
rect 545782 510938 545866 511174
rect 546102 510938 546134 511174
rect 545514 510854 546134 510938
rect 545514 510618 545546 510854
rect 545782 510618 545866 510854
rect 546102 510618 546134 510854
rect 545514 475174 546134 510618
rect 545514 474938 545546 475174
rect 545782 474938 545866 475174
rect 546102 474938 546134 475174
rect 545514 474854 546134 474938
rect 545514 474618 545546 474854
rect 545782 474618 545866 474854
rect 546102 474618 546134 474854
rect 545514 439174 546134 474618
rect 545514 438938 545546 439174
rect 545782 438938 545866 439174
rect 546102 438938 546134 439174
rect 545514 438854 546134 438938
rect 545514 438618 545546 438854
rect 545782 438618 545866 438854
rect 546102 438618 546134 438854
rect 545514 403174 546134 438618
rect 545514 402938 545546 403174
rect 545782 402938 545866 403174
rect 546102 402938 546134 403174
rect 545514 402854 546134 402938
rect 545514 402618 545546 402854
rect 545782 402618 545866 402854
rect 546102 402618 546134 402854
rect 545514 367174 546134 402618
rect 545514 366938 545546 367174
rect 545782 366938 545866 367174
rect 546102 366938 546134 367174
rect 545514 366854 546134 366938
rect 545514 366618 545546 366854
rect 545782 366618 545866 366854
rect 546102 366618 546134 366854
rect 545514 331174 546134 366618
rect 545514 330938 545546 331174
rect 545782 330938 545866 331174
rect 546102 330938 546134 331174
rect 545514 330854 546134 330938
rect 545514 330618 545546 330854
rect 545782 330618 545866 330854
rect 546102 330618 546134 330854
rect 545514 295174 546134 330618
rect 545514 294938 545546 295174
rect 545782 294938 545866 295174
rect 546102 294938 546134 295174
rect 545514 294854 546134 294938
rect 545514 294618 545546 294854
rect 545782 294618 545866 294854
rect 546102 294618 546134 294854
rect 545514 259174 546134 294618
rect 545514 258938 545546 259174
rect 545782 258938 545866 259174
rect 546102 258938 546134 259174
rect 545514 258854 546134 258938
rect 545514 258618 545546 258854
rect 545782 258618 545866 258854
rect 546102 258618 546134 258854
rect 545514 223174 546134 258618
rect 545514 222938 545546 223174
rect 545782 222938 545866 223174
rect 546102 222938 546134 223174
rect 545514 222854 546134 222938
rect 545514 222618 545546 222854
rect 545782 222618 545866 222854
rect 546102 222618 546134 222854
rect 545514 187174 546134 222618
rect 545514 186938 545546 187174
rect 545782 186938 545866 187174
rect 546102 186938 546134 187174
rect 545514 186854 546134 186938
rect 545514 186618 545546 186854
rect 545782 186618 545866 186854
rect 546102 186618 546134 186854
rect 545514 151174 546134 186618
rect 545514 150938 545546 151174
rect 545782 150938 545866 151174
rect 546102 150938 546134 151174
rect 545514 150854 546134 150938
rect 545514 150618 545546 150854
rect 545782 150618 545866 150854
rect 546102 150618 546134 150854
rect 545514 115174 546134 150618
rect 545514 114938 545546 115174
rect 545782 114938 545866 115174
rect 546102 114938 546134 115174
rect 545514 114854 546134 114938
rect 545514 114618 545546 114854
rect 545782 114618 545866 114854
rect 546102 114618 546134 114854
rect 545514 79174 546134 114618
rect 545514 78938 545546 79174
rect 545782 78938 545866 79174
rect 546102 78938 546134 79174
rect 545514 78854 546134 78938
rect 545514 78618 545546 78854
rect 545782 78618 545866 78854
rect 546102 78618 546134 78854
rect 545514 43174 546134 78618
rect 545514 42938 545546 43174
rect 545782 42938 545866 43174
rect 546102 42938 546134 43174
rect 545514 42854 546134 42938
rect 545514 42618 545546 42854
rect 545782 42618 545866 42854
rect 546102 42618 546134 42854
rect 545514 7174 546134 42618
rect 545514 6938 545546 7174
rect 545782 6938 545866 7174
rect 546102 6938 546134 7174
rect 545514 6854 546134 6938
rect 545514 6618 545546 6854
rect 545782 6618 545866 6854
rect 546102 6618 546134 6854
rect 545514 -2266 546134 6618
rect 545514 -2502 545546 -2266
rect 545782 -2502 545866 -2266
rect 546102 -2502 546134 -2266
rect 545514 -2586 546134 -2502
rect 545514 -2822 545546 -2586
rect 545782 -2822 545866 -2586
rect 546102 -2822 546134 -2586
rect 545514 -3814 546134 -2822
rect 549234 694894 549854 708122
rect 549234 694658 549266 694894
rect 549502 694658 549586 694894
rect 549822 694658 549854 694894
rect 549234 694574 549854 694658
rect 549234 694338 549266 694574
rect 549502 694338 549586 694574
rect 549822 694338 549854 694574
rect 549234 658894 549854 694338
rect 549234 658658 549266 658894
rect 549502 658658 549586 658894
rect 549822 658658 549854 658894
rect 549234 658574 549854 658658
rect 549234 658338 549266 658574
rect 549502 658338 549586 658574
rect 549822 658338 549854 658574
rect 549234 622894 549854 658338
rect 549234 622658 549266 622894
rect 549502 622658 549586 622894
rect 549822 622658 549854 622894
rect 549234 622574 549854 622658
rect 549234 622338 549266 622574
rect 549502 622338 549586 622574
rect 549822 622338 549854 622574
rect 549234 586894 549854 622338
rect 549234 586658 549266 586894
rect 549502 586658 549586 586894
rect 549822 586658 549854 586894
rect 549234 586574 549854 586658
rect 549234 586338 549266 586574
rect 549502 586338 549586 586574
rect 549822 586338 549854 586574
rect 549234 550894 549854 586338
rect 549234 550658 549266 550894
rect 549502 550658 549586 550894
rect 549822 550658 549854 550894
rect 549234 550574 549854 550658
rect 549234 550338 549266 550574
rect 549502 550338 549586 550574
rect 549822 550338 549854 550574
rect 549234 514894 549854 550338
rect 549234 514658 549266 514894
rect 549502 514658 549586 514894
rect 549822 514658 549854 514894
rect 549234 514574 549854 514658
rect 549234 514338 549266 514574
rect 549502 514338 549586 514574
rect 549822 514338 549854 514574
rect 549234 478894 549854 514338
rect 549234 478658 549266 478894
rect 549502 478658 549586 478894
rect 549822 478658 549854 478894
rect 549234 478574 549854 478658
rect 549234 478338 549266 478574
rect 549502 478338 549586 478574
rect 549822 478338 549854 478574
rect 549234 442894 549854 478338
rect 549234 442658 549266 442894
rect 549502 442658 549586 442894
rect 549822 442658 549854 442894
rect 549234 442574 549854 442658
rect 549234 442338 549266 442574
rect 549502 442338 549586 442574
rect 549822 442338 549854 442574
rect 549234 406894 549854 442338
rect 549234 406658 549266 406894
rect 549502 406658 549586 406894
rect 549822 406658 549854 406894
rect 549234 406574 549854 406658
rect 549234 406338 549266 406574
rect 549502 406338 549586 406574
rect 549822 406338 549854 406574
rect 549234 370894 549854 406338
rect 549234 370658 549266 370894
rect 549502 370658 549586 370894
rect 549822 370658 549854 370894
rect 549234 370574 549854 370658
rect 549234 370338 549266 370574
rect 549502 370338 549586 370574
rect 549822 370338 549854 370574
rect 549234 334894 549854 370338
rect 549234 334658 549266 334894
rect 549502 334658 549586 334894
rect 549822 334658 549854 334894
rect 549234 334574 549854 334658
rect 549234 334338 549266 334574
rect 549502 334338 549586 334574
rect 549822 334338 549854 334574
rect 549234 298894 549854 334338
rect 549234 298658 549266 298894
rect 549502 298658 549586 298894
rect 549822 298658 549854 298894
rect 549234 298574 549854 298658
rect 549234 298338 549266 298574
rect 549502 298338 549586 298574
rect 549822 298338 549854 298574
rect 549234 262894 549854 298338
rect 549234 262658 549266 262894
rect 549502 262658 549586 262894
rect 549822 262658 549854 262894
rect 549234 262574 549854 262658
rect 549234 262338 549266 262574
rect 549502 262338 549586 262574
rect 549822 262338 549854 262574
rect 549234 226894 549854 262338
rect 549234 226658 549266 226894
rect 549502 226658 549586 226894
rect 549822 226658 549854 226894
rect 549234 226574 549854 226658
rect 549234 226338 549266 226574
rect 549502 226338 549586 226574
rect 549822 226338 549854 226574
rect 549234 190894 549854 226338
rect 549234 190658 549266 190894
rect 549502 190658 549586 190894
rect 549822 190658 549854 190894
rect 549234 190574 549854 190658
rect 549234 190338 549266 190574
rect 549502 190338 549586 190574
rect 549822 190338 549854 190574
rect 549234 154894 549854 190338
rect 549234 154658 549266 154894
rect 549502 154658 549586 154894
rect 549822 154658 549854 154894
rect 549234 154574 549854 154658
rect 549234 154338 549266 154574
rect 549502 154338 549586 154574
rect 549822 154338 549854 154574
rect 549234 118894 549854 154338
rect 549234 118658 549266 118894
rect 549502 118658 549586 118894
rect 549822 118658 549854 118894
rect 549234 118574 549854 118658
rect 549234 118338 549266 118574
rect 549502 118338 549586 118574
rect 549822 118338 549854 118574
rect 549234 82894 549854 118338
rect 549234 82658 549266 82894
rect 549502 82658 549586 82894
rect 549822 82658 549854 82894
rect 549234 82574 549854 82658
rect 549234 82338 549266 82574
rect 549502 82338 549586 82574
rect 549822 82338 549854 82574
rect 549234 46894 549854 82338
rect 549234 46658 549266 46894
rect 549502 46658 549586 46894
rect 549822 46658 549854 46894
rect 549234 46574 549854 46658
rect 549234 46338 549266 46574
rect 549502 46338 549586 46574
rect 549822 46338 549854 46574
rect 549234 10894 549854 46338
rect 549234 10658 549266 10894
rect 549502 10658 549586 10894
rect 549822 10658 549854 10894
rect 549234 10574 549854 10658
rect 549234 10338 549266 10574
rect 549502 10338 549586 10574
rect 549822 10338 549854 10574
rect 549234 -4186 549854 10338
rect 549234 -4422 549266 -4186
rect 549502 -4422 549586 -4186
rect 549822 -4422 549854 -4186
rect 549234 -4506 549854 -4422
rect 549234 -4742 549266 -4506
rect 549502 -4742 549586 -4506
rect 549822 -4742 549854 -4506
rect 549234 -5734 549854 -4742
rect 552954 698614 553574 710042
rect 570954 711558 571574 711590
rect 570954 711322 570986 711558
rect 571222 711322 571306 711558
rect 571542 711322 571574 711558
rect 570954 711238 571574 711322
rect 570954 711002 570986 711238
rect 571222 711002 571306 711238
rect 571542 711002 571574 711238
rect 567234 709638 567854 709670
rect 567234 709402 567266 709638
rect 567502 709402 567586 709638
rect 567822 709402 567854 709638
rect 567234 709318 567854 709402
rect 567234 709082 567266 709318
rect 567502 709082 567586 709318
rect 567822 709082 567854 709318
rect 563514 707718 564134 707750
rect 563514 707482 563546 707718
rect 563782 707482 563866 707718
rect 564102 707482 564134 707718
rect 563514 707398 564134 707482
rect 563514 707162 563546 707398
rect 563782 707162 563866 707398
rect 564102 707162 564134 707398
rect 552954 698378 552986 698614
rect 553222 698378 553306 698614
rect 553542 698378 553574 698614
rect 552954 698294 553574 698378
rect 552954 698058 552986 698294
rect 553222 698058 553306 698294
rect 553542 698058 553574 698294
rect 552954 662614 553574 698058
rect 552954 662378 552986 662614
rect 553222 662378 553306 662614
rect 553542 662378 553574 662614
rect 552954 662294 553574 662378
rect 552954 662058 552986 662294
rect 553222 662058 553306 662294
rect 553542 662058 553574 662294
rect 552954 626614 553574 662058
rect 552954 626378 552986 626614
rect 553222 626378 553306 626614
rect 553542 626378 553574 626614
rect 552954 626294 553574 626378
rect 552954 626058 552986 626294
rect 553222 626058 553306 626294
rect 553542 626058 553574 626294
rect 552954 590614 553574 626058
rect 552954 590378 552986 590614
rect 553222 590378 553306 590614
rect 553542 590378 553574 590614
rect 552954 590294 553574 590378
rect 552954 590058 552986 590294
rect 553222 590058 553306 590294
rect 553542 590058 553574 590294
rect 552954 554614 553574 590058
rect 552954 554378 552986 554614
rect 553222 554378 553306 554614
rect 553542 554378 553574 554614
rect 552954 554294 553574 554378
rect 552954 554058 552986 554294
rect 553222 554058 553306 554294
rect 553542 554058 553574 554294
rect 552954 518614 553574 554058
rect 552954 518378 552986 518614
rect 553222 518378 553306 518614
rect 553542 518378 553574 518614
rect 552954 518294 553574 518378
rect 552954 518058 552986 518294
rect 553222 518058 553306 518294
rect 553542 518058 553574 518294
rect 552954 482614 553574 518058
rect 552954 482378 552986 482614
rect 553222 482378 553306 482614
rect 553542 482378 553574 482614
rect 552954 482294 553574 482378
rect 552954 482058 552986 482294
rect 553222 482058 553306 482294
rect 553542 482058 553574 482294
rect 552954 446614 553574 482058
rect 552954 446378 552986 446614
rect 553222 446378 553306 446614
rect 553542 446378 553574 446614
rect 552954 446294 553574 446378
rect 552954 446058 552986 446294
rect 553222 446058 553306 446294
rect 553542 446058 553574 446294
rect 552954 410614 553574 446058
rect 552954 410378 552986 410614
rect 553222 410378 553306 410614
rect 553542 410378 553574 410614
rect 552954 410294 553574 410378
rect 552954 410058 552986 410294
rect 553222 410058 553306 410294
rect 553542 410058 553574 410294
rect 552954 374614 553574 410058
rect 552954 374378 552986 374614
rect 553222 374378 553306 374614
rect 553542 374378 553574 374614
rect 552954 374294 553574 374378
rect 552954 374058 552986 374294
rect 553222 374058 553306 374294
rect 553542 374058 553574 374294
rect 552954 338614 553574 374058
rect 552954 338378 552986 338614
rect 553222 338378 553306 338614
rect 553542 338378 553574 338614
rect 552954 338294 553574 338378
rect 552954 338058 552986 338294
rect 553222 338058 553306 338294
rect 553542 338058 553574 338294
rect 552954 302614 553574 338058
rect 552954 302378 552986 302614
rect 553222 302378 553306 302614
rect 553542 302378 553574 302614
rect 552954 302294 553574 302378
rect 552954 302058 552986 302294
rect 553222 302058 553306 302294
rect 553542 302058 553574 302294
rect 552954 266614 553574 302058
rect 552954 266378 552986 266614
rect 553222 266378 553306 266614
rect 553542 266378 553574 266614
rect 552954 266294 553574 266378
rect 552954 266058 552986 266294
rect 553222 266058 553306 266294
rect 553542 266058 553574 266294
rect 552954 230614 553574 266058
rect 552954 230378 552986 230614
rect 553222 230378 553306 230614
rect 553542 230378 553574 230614
rect 552954 230294 553574 230378
rect 552954 230058 552986 230294
rect 553222 230058 553306 230294
rect 553542 230058 553574 230294
rect 552954 194614 553574 230058
rect 552954 194378 552986 194614
rect 553222 194378 553306 194614
rect 553542 194378 553574 194614
rect 552954 194294 553574 194378
rect 552954 194058 552986 194294
rect 553222 194058 553306 194294
rect 553542 194058 553574 194294
rect 552954 158614 553574 194058
rect 552954 158378 552986 158614
rect 553222 158378 553306 158614
rect 553542 158378 553574 158614
rect 552954 158294 553574 158378
rect 552954 158058 552986 158294
rect 553222 158058 553306 158294
rect 553542 158058 553574 158294
rect 552954 122614 553574 158058
rect 552954 122378 552986 122614
rect 553222 122378 553306 122614
rect 553542 122378 553574 122614
rect 552954 122294 553574 122378
rect 552954 122058 552986 122294
rect 553222 122058 553306 122294
rect 553542 122058 553574 122294
rect 552954 86614 553574 122058
rect 552954 86378 552986 86614
rect 553222 86378 553306 86614
rect 553542 86378 553574 86614
rect 552954 86294 553574 86378
rect 552954 86058 552986 86294
rect 553222 86058 553306 86294
rect 553542 86058 553574 86294
rect 552954 50614 553574 86058
rect 552954 50378 552986 50614
rect 553222 50378 553306 50614
rect 553542 50378 553574 50614
rect 552954 50294 553574 50378
rect 552954 50058 552986 50294
rect 553222 50058 553306 50294
rect 553542 50058 553574 50294
rect 552954 14614 553574 50058
rect 552954 14378 552986 14614
rect 553222 14378 553306 14614
rect 553542 14378 553574 14614
rect 552954 14294 553574 14378
rect 552954 14058 552986 14294
rect 553222 14058 553306 14294
rect 553542 14058 553574 14294
rect 534954 -7302 534986 -7066
rect 535222 -7302 535306 -7066
rect 535542 -7302 535574 -7066
rect 534954 -7386 535574 -7302
rect 534954 -7622 534986 -7386
rect 535222 -7622 535306 -7386
rect 535542 -7622 535574 -7386
rect 534954 -7654 535574 -7622
rect 552954 -6106 553574 14058
rect 559794 705798 560414 705830
rect 559794 705562 559826 705798
rect 560062 705562 560146 705798
rect 560382 705562 560414 705798
rect 559794 705478 560414 705562
rect 559794 705242 559826 705478
rect 560062 705242 560146 705478
rect 560382 705242 560414 705478
rect 559794 669454 560414 705242
rect 559794 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 560414 669454
rect 559794 669134 560414 669218
rect 559794 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 560414 669134
rect 559794 633454 560414 668898
rect 559794 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 560414 633454
rect 559794 633134 560414 633218
rect 559794 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 560414 633134
rect 559794 597454 560414 632898
rect 559794 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 560414 597454
rect 559794 597134 560414 597218
rect 559794 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 560414 597134
rect 559794 561454 560414 596898
rect 559794 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 560414 561454
rect 559794 561134 560414 561218
rect 559794 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 560414 561134
rect 559794 525454 560414 560898
rect 559794 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 560414 525454
rect 559794 525134 560414 525218
rect 559794 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 560414 525134
rect 559794 489454 560414 524898
rect 559794 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 560414 489454
rect 559794 489134 560414 489218
rect 559794 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 560414 489134
rect 559794 453454 560414 488898
rect 559794 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 560414 453454
rect 559794 453134 560414 453218
rect 559794 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 560414 453134
rect 559794 417454 560414 452898
rect 559794 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 560414 417454
rect 559794 417134 560414 417218
rect 559794 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 560414 417134
rect 559794 381454 560414 416898
rect 559794 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 560414 381454
rect 559794 381134 560414 381218
rect 559794 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 560414 381134
rect 559794 345454 560414 380898
rect 559794 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 560414 345454
rect 559794 345134 560414 345218
rect 559794 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 560414 345134
rect 559794 309454 560414 344898
rect 559794 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 560414 309454
rect 559794 309134 560414 309218
rect 559794 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 560414 309134
rect 559794 273454 560414 308898
rect 559794 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 560414 273454
rect 559794 273134 560414 273218
rect 559794 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 560414 273134
rect 559794 237454 560414 272898
rect 559794 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 560414 237454
rect 559794 237134 560414 237218
rect 559794 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 560414 237134
rect 559794 201454 560414 236898
rect 559794 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 560414 201454
rect 559794 201134 560414 201218
rect 559794 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 560414 201134
rect 559794 165454 560414 200898
rect 559794 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 560414 165454
rect 559794 165134 560414 165218
rect 559794 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 560414 165134
rect 559794 129454 560414 164898
rect 559794 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 560414 129454
rect 559794 129134 560414 129218
rect 559794 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 560414 129134
rect 559794 93454 560414 128898
rect 559794 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 560414 93454
rect 559794 93134 560414 93218
rect 559794 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 560414 93134
rect 559794 57454 560414 92898
rect 559794 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 560414 57454
rect 559794 57134 560414 57218
rect 559794 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 560414 57134
rect 559794 21454 560414 56898
rect 559794 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 560414 21454
rect 559794 21134 560414 21218
rect 559794 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 560414 21134
rect 559794 -1306 560414 20898
rect 559794 -1542 559826 -1306
rect 560062 -1542 560146 -1306
rect 560382 -1542 560414 -1306
rect 559794 -1626 560414 -1542
rect 559794 -1862 559826 -1626
rect 560062 -1862 560146 -1626
rect 560382 -1862 560414 -1626
rect 559794 -1894 560414 -1862
rect 563514 673174 564134 707162
rect 563514 672938 563546 673174
rect 563782 672938 563866 673174
rect 564102 672938 564134 673174
rect 563514 672854 564134 672938
rect 563514 672618 563546 672854
rect 563782 672618 563866 672854
rect 564102 672618 564134 672854
rect 563514 637174 564134 672618
rect 563514 636938 563546 637174
rect 563782 636938 563866 637174
rect 564102 636938 564134 637174
rect 563514 636854 564134 636938
rect 563514 636618 563546 636854
rect 563782 636618 563866 636854
rect 564102 636618 564134 636854
rect 563514 601174 564134 636618
rect 563514 600938 563546 601174
rect 563782 600938 563866 601174
rect 564102 600938 564134 601174
rect 563514 600854 564134 600938
rect 563514 600618 563546 600854
rect 563782 600618 563866 600854
rect 564102 600618 564134 600854
rect 563514 565174 564134 600618
rect 563514 564938 563546 565174
rect 563782 564938 563866 565174
rect 564102 564938 564134 565174
rect 563514 564854 564134 564938
rect 563514 564618 563546 564854
rect 563782 564618 563866 564854
rect 564102 564618 564134 564854
rect 563514 529174 564134 564618
rect 563514 528938 563546 529174
rect 563782 528938 563866 529174
rect 564102 528938 564134 529174
rect 563514 528854 564134 528938
rect 563514 528618 563546 528854
rect 563782 528618 563866 528854
rect 564102 528618 564134 528854
rect 563514 493174 564134 528618
rect 563514 492938 563546 493174
rect 563782 492938 563866 493174
rect 564102 492938 564134 493174
rect 563514 492854 564134 492938
rect 563514 492618 563546 492854
rect 563782 492618 563866 492854
rect 564102 492618 564134 492854
rect 563514 457174 564134 492618
rect 563514 456938 563546 457174
rect 563782 456938 563866 457174
rect 564102 456938 564134 457174
rect 563514 456854 564134 456938
rect 563514 456618 563546 456854
rect 563782 456618 563866 456854
rect 564102 456618 564134 456854
rect 563514 421174 564134 456618
rect 563514 420938 563546 421174
rect 563782 420938 563866 421174
rect 564102 420938 564134 421174
rect 563514 420854 564134 420938
rect 563514 420618 563546 420854
rect 563782 420618 563866 420854
rect 564102 420618 564134 420854
rect 563514 385174 564134 420618
rect 563514 384938 563546 385174
rect 563782 384938 563866 385174
rect 564102 384938 564134 385174
rect 563514 384854 564134 384938
rect 563514 384618 563546 384854
rect 563782 384618 563866 384854
rect 564102 384618 564134 384854
rect 563514 349174 564134 384618
rect 563514 348938 563546 349174
rect 563782 348938 563866 349174
rect 564102 348938 564134 349174
rect 563514 348854 564134 348938
rect 563514 348618 563546 348854
rect 563782 348618 563866 348854
rect 564102 348618 564134 348854
rect 563514 313174 564134 348618
rect 563514 312938 563546 313174
rect 563782 312938 563866 313174
rect 564102 312938 564134 313174
rect 563514 312854 564134 312938
rect 563514 312618 563546 312854
rect 563782 312618 563866 312854
rect 564102 312618 564134 312854
rect 563514 277174 564134 312618
rect 563514 276938 563546 277174
rect 563782 276938 563866 277174
rect 564102 276938 564134 277174
rect 563514 276854 564134 276938
rect 563514 276618 563546 276854
rect 563782 276618 563866 276854
rect 564102 276618 564134 276854
rect 563514 241174 564134 276618
rect 563514 240938 563546 241174
rect 563782 240938 563866 241174
rect 564102 240938 564134 241174
rect 563514 240854 564134 240938
rect 563514 240618 563546 240854
rect 563782 240618 563866 240854
rect 564102 240618 564134 240854
rect 563514 205174 564134 240618
rect 563514 204938 563546 205174
rect 563782 204938 563866 205174
rect 564102 204938 564134 205174
rect 563514 204854 564134 204938
rect 563514 204618 563546 204854
rect 563782 204618 563866 204854
rect 564102 204618 564134 204854
rect 563514 169174 564134 204618
rect 563514 168938 563546 169174
rect 563782 168938 563866 169174
rect 564102 168938 564134 169174
rect 563514 168854 564134 168938
rect 563514 168618 563546 168854
rect 563782 168618 563866 168854
rect 564102 168618 564134 168854
rect 563514 133174 564134 168618
rect 563514 132938 563546 133174
rect 563782 132938 563866 133174
rect 564102 132938 564134 133174
rect 563514 132854 564134 132938
rect 563514 132618 563546 132854
rect 563782 132618 563866 132854
rect 564102 132618 564134 132854
rect 563514 97174 564134 132618
rect 563514 96938 563546 97174
rect 563782 96938 563866 97174
rect 564102 96938 564134 97174
rect 563514 96854 564134 96938
rect 563514 96618 563546 96854
rect 563782 96618 563866 96854
rect 564102 96618 564134 96854
rect 563514 61174 564134 96618
rect 563514 60938 563546 61174
rect 563782 60938 563866 61174
rect 564102 60938 564134 61174
rect 563514 60854 564134 60938
rect 563514 60618 563546 60854
rect 563782 60618 563866 60854
rect 564102 60618 564134 60854
rect 563514 25174 564134 60618
rect 563514 24938 563546 25174
rect 563782 24938 563866 25174
rect 564102 24938 564134 25174
rect 563514 24854 564134 24938
rect 563514 24618 563546 24854
rect 563782 24618 563866 24854
rect 564102 24618 564134 24854
rect 563514 -3226 564134 24618
rect 563514 -3462 563546 -3226
rect 563782 -3462 563866 -3226
rect 564102 -3462 564134 -3226
rect 563514 -3546 564134 -3462
rect 563514 -3782 563546 -3546
rect 563782 -3782 563866 -3546
rect 564102 -3782 564134 -3546
rect 563514 -3814 564134 -3782
rect 567234 676894 567854 709082
rect 567234 676658 567266 676894
rect 567502 676658 567586 676894
rect 567822 676658 567854 676894
rect 567234 676574 567854 676658
rect 567234 676338 567266 676574
rect 567502 676338 567586 676574
rect 567822 676338 567854 676574
rect 567234 640894 567854 676338
rect 567234 640658 567266 640894
rect 567502 640658 567586 640894
rect 567822 640658 567854 640894
rect 567234 640574 567854 640658
rect 567234 640338 567266 640574
rect 567502 640338 567586 640574
rect 567822 640338 567854 640574
rect 567234 604894 567854 640338
rect 567234 604658 567266 604894
rect 567502 604658 567586 604894
rect 567822 604658 567854 604894
rect 567234 604574 567854 604658
rect 567234 604338 567266 604574
rect 567502 604338 567586 604574
rect 567822 604338 567854 604574
rect 567234 568894 567854 604338
rect 567234 568658 567266 568894
rect 567502 568658 567586 568894
rect 567822 568658 567854 568894
rect 567234 568574 567854 568658
rect 567234 568338 567266 568574
rect 567502 568338 567586 568574
rect 567822 568338 567854 568574
rect 567234 532894 567854 568338
rect 567234 532658 567266 532894
rect 567502 532658 567586 532894
rect 567822 532658 567854 532894
rect 567234 532574 567854 532658
rect 567234 532338 567266 532574
rect 567502 532338 567586 532574
rect 567822 532338 567854 532574
rect 567234 496894 567854 532338
rect 567234 496658 567266 496894
rect 567502 496658 567586 496894
rect 567822 496658 567854 496894
rect 567234 496574 567854 496658
rect 567234 496338 567266 496574
rect 567502 496338 567586 496574
rect 567822 496338 567854 496574
rect 567234 460894 567854 496338
rect 567234 460658 567266 460894
rect 567502 460658 567586 460894
rect 567822 460658 567854 460894
rect 567234 460574 567854 460658
rect 567234 460338 567266 460574
rect 567502 460338 567586 460574
rect 567822 460338 567854 460574
rect 567234 424894 567854 460338
rect 567234 424658 567266 424894
rect 567502 424658 567586 424894
rect 567822 424658 567854 424894
rect 567234 424574 567854 424658
rect 567234 424338 567266 424574
rect 567502 424338 567586 424574
rect 567822 424338 567854 424574
rect 567234 388894 567854 424338
rect 567234 388658 567266 388894
rect 567502 388658 567586 388894
rect 567822 388658 567854 388894
rect 567234 388574 567854 388658
rect 567234 388338 567266 388574
rect 567502 388338 567586 388574
rect 567822 388338 567854 388574
rect 567234 352894 567854 388338
rect 567234 352658 567266 352894
rect 567502 352658 567586 352894
rect 567822 352658 567854 352894
rect 567234 352574 567854 352658
rect 567234 352338 567266 352574
rect 567502 352338 567586 352574
rect 567822 352338 567854 352574
rect 567234 316894 567854 352338
rect 567234 316658 567266 316894
rect 567502 316658 567586 316894
rect 567822 316658 567854 316894
rect 567234 316574 567854 316658
rect 567234 316338 567266 316574
rect 567502 316338 567586 316574
rect 567822 316338 567854 316574
rect 567234 280894 567854 316338
rect 567234 280658 567266 280894
rect 567502 280658 567586 280894
rect 567822 280658 567854 280894
rect 567234 280574 567854 280658
rect 567234 280338 567266 280574
rect 567502 280338 567586 280574
rect 567822 280338 567854 280574
rect 567234 244894 567854 280338
rect 567234 244658 567266 244894
rect 567502 244658 567586 244894
rect 567822 244658 567854 244894
rect 567234 244574 567854 244658
rect 567234 244338 567266 244574
rect 567502 244338 567586 244574
rect 567822 244338 567854 244574
rect 567234 208894 567854 244338
rect 567234 208658 567266 208894
rect 567502 208658 567586 208894
rect 567822 208658 567854 208894
rect 567234 208574 567854 208658
rect 567234 208338 567266 208574
rect 567502 208338 567586 208574
rect 567822 208338 567854 208574
rect 567234 172894 567854 208338
rect 567234 172658 567266 172894
rect 567502 172658 567586 172894
rect 567822 172658 567854 172894
rect 567234 172574 567854 172658
rect 567234 172338 567266 172574
rect 567502 172338 567586 172574
rect 567822 172338 567854 172574
rect 567234 136894 567854 172338
rect 567234 136658 567266 136894
rect 567502 136658 567586 136894
rect 567822 136658 567854 136894
rect 567234 136574 567854 136658
rect 567234 136338 567266 136574
rect 567502 136338 567586 136574
rect 567822 136338 567854 136574
rect 567234 100894 567854 136338
rect 567234 100658 567266 100894
rect 567502 100658 567586 100894
rect 567822 100658 567854 100894
rect 567234 100574 567854 100658
rect 567234 100338 567266 100574
rect 567502 100338 567586 100574
rect 567822 100338 567854 100574
rect 567234 64894 567854 100338
rect 567234 64658 567266 64894
rect 567502 64658 567586 64894
rect 567822 64658 567854 64894
rect 567234 64574 567854 64658
rect 567234 64338 567266 64574
rect 567502 64338 567586 64574
rect 567822 64338 567854 64574
rect 567234 28894 567854 64338
rect 567234 28658 567266 28894
rect 567502 28658 567586 28894
rect 567822 28658 567854 28894
rect 567234 28574 567854 28658
rect 567234 28338 567266 28574
rect 567502 28338 567586 28574
rect 567822 28338 567854 28574
rect 567234 -5146 567854 28338
rect 567234 -5382 567266 -5146
rect 567502 -5382 567586 -5146
rect 567822 -5382 567854 -5146
rect 567234 -5466 567854 -5382
rect 567234 -5702 567266 -5466
rect 567502 -5702 567586 -5466
rect 567822 -5702 567854 -5466
rect 567234 -5734 567854 -5702
rect 570954 680614 571574 711002
rect 592030 711558 592650 711590
rect 592030 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect 592030 711238 592650 711322
rect 592030 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect 591070 710598 591690 710630
rect 591070 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect 591070 710278 591690 710362
rect 591070 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect 590110 709638 590730 709670
rect 590110 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect 590110 709318 590730 709402
rect 590110 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect 589150 708678 589770 708710
rect 589150 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect 589150 708358 589770 708442
rect 589150 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect 581514 706758 582134 707750
rect 588190 707718 588810 707750
rect 588190 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect 588190 707398 588810 707482
rect 588190 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect 581514 706522 581546 706758
rect 581782 706522 581866 706758
rect 582102 706522 582134 706758
rect 581514 706438 582134 706522
rect 581514 706202 581546 706438
rect 581782 706202 581866 706438
rect 582102 706202 582134 706438
rect 570954 680378 570986 680614
rect 571222 680378 571306 680614
rect 571542 680378 571574 680614
rect 570954 680294 571574 680378
rect 570954 680058 570986 680294
rect 571222 680058 571306 680294
rect 571542 680058 571574 680294
rect 570954 644614 571574 680058
rect 570954 644378 570986 644614
rect 571222 644378 571306 644614
rect 571542 644378 571574 644614
rect 570954 644294 571574 644378
rect 570954 644058 570986 644294
rect 571222 644058 571306 644294
rect 571542 644058 571574 644294
rect 570954 608614 571574 644058
rect 570954 608378 570986 608614
rect 571222 608378 571306 608614
rect 571542 608378 571574 608614
rect 570954 608294 571574 608378
rect 570954 608058 570986 608294
rect 571222 608058 571306 608294
rect 571542 608058 571574 608294
rect 570954 572614 571574 608058
rect 570954 572378 570986 572614
rect 571222 572378 571306 572614
rect 571542 572378 571574 572614
rect 570954 572294 571574 572378
rect 570954 572058 570986 572294
rect 571222 572058 571306 572294
rect 571542 572058 571574 572294
rect 570954 536614 571574 572058
rect 570954 536378 570986 536614
rect 571222 536378 571306 536614
rect 571542 536378 571574 536614
rect 570954 536294 571574 536378
rect 570954 536058 570986 536294
rect 571222 536058 571306 536294
rect 571542 536058 571574 536294
rect 570954 500614 571574 536058
rect 570954 500378 570986 500614
rect 571222 500378 571306 500614
rect 571542 500378 571574 500614
rect 570954 500294 571574 500378
rect 570954 500058 570986 500294
rect 571222 500058 571306 500294
rect 571542 500058 571574 500294
rect 570954 464614 571574 500058
rect 570954 464378 570986 464614
rect 571222 464378 571306 464614
rect 571542 464378 571574 464614
rect 570954 464294 571574 464378
rect 570954 464058 570986 464294
rect 571222 464058 571306 464294
rect 571542 464058 571574 464294
rect 570954 428614 571574 464058
rect 570954 428378 570986 428614
rect 571222 428378 571306 428614
rect 571542 428378 571574 428614
rect 570954 428294 571574 428378
rect 570954 428058 570986 428294
rect 571222 428058 571306 428294
rect 571542 428058 571574 428294
rect 570954 392614 571574 428058
rect 570954 392378 570986 392614
rect 571222 392378 571306 392614
rect 571542 392378 571574 392614
rect 570954 392294 571574 392378
rect 570954 392058 570986 392294
rect 571222 392058 571306 392294
rect 571542 392058 571574 392294
rect 570954 356614 571574 392058
rect 570954 356378 570986 356614
rect 571222 356378 571306 356614
rect 571542 356378 571574 356614
rect 570954 356294 571574 356378
rect 570954 356058 570986 356294
rect 571222 356058 571306 356294
rect 571542 356058 571574 356294
rect 570954 320614 571574 356058
rect 570954 320378 570986 320614
rect 571222 320378 571306 320614
rect 571542 320378 571574 320614
rect 570954 320294 571574 320378
rect 570954 320058 570986 320294
rect 571222 320058 571306 320294
rect 571542 320058 571574 320294
rect 570954 284614 571574 320058
rect 570954 284378 570986 284614
rect 571222 284378 571306 284614
rect 571542 284378 571574 284614
rect 570954 284294 571574 284378
rect 570954 284058 570986 284294
rect 571222 284058 571306 284294
rect 571542 284058 571574 284294
rect 570954 248614 571574 284058
rect 570954 248378 570986 248614
rect 571222 248378 571306 248614
rect 571542 248378 571574 248614
rect 570954 248294 571574 248378
rect 570954 248058 570986 248294
rect 571222 248058 571306 248294
rect 571542 248058 571574 248294
rect 570954 212614 571574 248058
rect 570954 212378 570986 212614
rect 571222 212378 571306 212614
rect 571542 212378 571574 212614
rect 570954 212294 571574 212378
rect 570954 212058 570986 212294
rect 571222 212058 571306 212294
rect 571542 212058 571574 212294
rect 570954 176614 571574 212058
rect 570954 176378 570986 176614
rect 571222 176378 571306 176614
rect 571542 176378 571574 176614
rect 570954 176294 571574 176378
rect 570954 176058 570986 176294
rect 571222 176058 571306 176294
rect 571542 176058 571574 176294
rect 570954 140614 571574 176058
rect 570954 140378 570986 140614
rect 571222 140378 571306 140614
rect 571542 140378 571574 140614
rect 570954 140294 571574 140378
rect 570954 140058 570986 140294
rect 571222 140058 571306 140294
rect 571542 140058 571574 140294
rect 570954 104614 571574 140058
rect 570954 104378 570986 104614
rect 571222 104378 571306 104614
rect 571542 104378 571574 104614
rect 570954 104294 571574 104378
rect 570954 104058 570986 104294
rect 571222 104058 571306 104294
rect 571542 104058 571574 104294
rect 570954 68614 571574 104058
rect 570954 68378 570986 68614
rect 571222 68378 571306 68614
rect 571542 68378 571574 68614
rect 570954 68294 571574 68378
rect 570954 68058 570986 68294
rect 571222 68058 571306 68294
rect 571542 68058 571574 68294
rect 570954 32614 571574 68058
rect 570954 32378 570986 32614
rect 571222 32378 571306 32614
rect 571542 32378 571574 32614
rect 570954 32294 571574 32378
rect 570954 32058 570986 32294
rect 571222 32058 571306 32294
rect 571542 32058 571574 32294
rect 552954 -6342 552986 -6106
rect 553222 -6342 553306 -6106
rect 553542 -6342 553574 -6106
rect 552954 -6426 553574 -6342
rect 552954 -6662 552986 -6426
rect 553222 -6662 553306 -6426
rect 553542 -6662 553574 -6426
rect 552954 -7654 553574 -6662
rect 570954 -7066 571574 32058
rect 577794 704838 578414 705830
rect 577794 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 578414 704838
rect 577794 704518 578414 704602
rect 577794 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 578414 704518
rect 577794 687454 578414 704282
rect 577794 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 578414 687454
rect 577794 687134 578414 687218
rect 577794 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 578414 687134
rect 577794 651454 578414 686898
rect 577794 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 578414 651454
rect 577794 651134 578414 651218
rect 577794 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 578414 651134
rect 577794 615454 578414 650898
rect 577794 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 578414 615454
rect 577794 615134 578414 615218
rect 577794 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 578414 615134
rect 577794 579454 578414 614898
rect 577794 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 578414 579454
rect 577794 579134 578414 579218
rect 577794 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 578414 579134
rect 577794 543454 578414 578898
rect 577794 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 578414 543454
rect 577794 543134 578414 543218
rect 577794 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 578414 543134
rect 577794 507454 578414 542898
rect 577794 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 578414 507454
rect 577794 507134 578414 507218
rect 577794 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 578414 507134
rect 577794 471454 578414 506898
rect 577794 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 578414 471454
rect 577794 471134 578414 471218
rect 577794 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 578414 471134
rect 577794 435454 578414 470898
rect 577794 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 578414 435454
rect 577794 435134 578414 435218
rect 577794 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 578414 435134
rect 577794 399454 578414 434898
rect 577794 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 578414 399454
rect 577794 399134 578414 399218
rect 577794 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 578414 399134
rect 577794 363454 578414 398898
rect 577794 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 578414 363454
rect 577794 363134 578414 363218
rect 577794 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 578414 363134
rect 577794 327454 578414 362898
rect 577794 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 578414 327454
rect 577794 327134 578414 327218
rect 577794 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 578414 327134
rect 577794 291454 578414 326898
rect 577794 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 578414 291454
rect 577794 291134 578414 291218
rect 577794 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 578414 291134
rect 577794 255454 578414 290898
rect 577794 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 578414 255454
rect 577794 255134 578414 255218
rect 577794 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 578414 255134
rect 577794 219454 578414 254898
rect 577794 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 578414 219454
rect 577794 219134 578414 219218
rect 577794 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 578414 219134
rect 577794 183454 578414 218898
rect 577794 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 578414 183454
rect 577794 183134 578414 183218
rect 577794 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 578414 183134
rect 577794 147454 578414 182898
rect 577794 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 578414 147454
rect 577794 147134 578414 147218
rect 577794 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 578414 147134
rect 577794 111454 578414 146898
rect 577794 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 578414 111454
rect 577794 111134 578414 111218
rect 577794 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 578414 111134
rect 577794 75454 578414 110898
rect 577794 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 578414 75454
rect 577794 75134 578414 75218
rect 577794 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 578414 75134
rect 577794 39454 578414 74898
rect 577794 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 578414 39454
rect 577794 39134 578414 39218
rect 577794 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 578414 39134
rect 577794 3454 578414 38898
rect 577794 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 578414 3454
rect 577794 3134 578414 3218
rect 577794 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 578414 3134
rect 577794 -346 578414 2898
rect 577794 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 578414 -346
rect 577794 -666 578414 -582
rect 577794 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 578414 -666
rect 577794 -1894 578414 -902
rect 581514 691174 582134 706202
rect 587230 706758 587850 706790
rect 587230 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect 587230 706438 587850 706522
rect 587230 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect 586270 705798 586890 705830
rect 586270 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect 586270 705478 586890 705562
rect 586270 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect 581514 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 582134 691174
rect 581514 690854 582134 690938
rect 581514 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 582134 690854
rect 581514 655174 582134 690618
rect 581514 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 582134 655174
rect 581514 654854 582134 654938
rect 581514 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 582134 654854
rect 581514 619174 582134 654618
rect 581514 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 582134 619174
rect 581514 618854 582134 618938
rect 581514 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 582134 618854
rect 581514 583174 582134 618618
rect 581514 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 582134 583174
rect 581514 582854 582134 582938
rect 581514 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 582134 582854
rect 581514 547174 582134 582618
rect 581514 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 582134 547174
rect 581514 546854 582134 546938
rect 581514 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 582134 546854
rect 581514 511174 582134 546618
rect 581514 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 582134 511174
rect 581514 510854 582134 510938
rect 581514 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 582134 510854
rect 581514 475174 582134 510618
rect 581514 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 582134 475174
rect 581514 474854 582134 474938
rect 581514 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 582134 474854
rect 581514 439174 582134 474618
rect 581514 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 582134 439174
rect 581514 438854 582134 438938
rect 581514 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 582134 438854
rect 581514 403174 582134 438618
rect 581514 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 582134 403174
rect 581514 402854 582134 402938
rect 581514 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 582134 402854
rect 581514 367174 582134 402618
rect 581514 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 582134 367174
rect 581514 366854 582134 366938
rect 581514 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 582134 366854
rect 581514 331174 582134 366618
rect 581514 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 582134 331174
rect 581514 330854 582134 330938
rect 581514 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 582134 330854
rect 581514 295174 582134 330618
rect 581514 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 582134 295174
rect 581514 294854 582134 294938
rect 581514 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 582134 294854
rect 581514 259174 582134 294618
rect 581514 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 582134 259174
rect 581514 258854 582134 258938
rect 581514 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 582134 258854
rect 581514 223174 582134 258618
rect 581514 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 582134 223174
rect 581514 222854 582134 222938
rect 581514 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 582134 222854
rect 581514 187174 582134 222618
rect 581514 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 582134 187174
rect 581514 186854 582134 186938
rect 581514 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 582134 186854
rect 581514 151174 582134 186618
rect 581514 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 582134 151174
rect 581514 150854 582134 150938
rect 581514 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 582134 150854
rect 581514 115174 582134 150618
rect 581514 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 582134 115174
rect 581514 114854 582134 114938
rect 581514 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 582134 114854
rect 581514 79174 582134 114618
rect 581514 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 582134 79174
rect 581514 78854 582134 78938
rect 581514 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 582134 78854
rect 581514 43174 582134 78618
rect 581514 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 582134 43174
rect 581514 42854 582134 42938
rect 581514 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 582134 42854
rect 581514 7174 582134 42618
rect 581514 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 582134 7174
rect 581514 6854 582134 6938
rect 581514 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 582134 6854
rect 581514 -2266 582134 6618
rect 585310 704838 585930 704870
rect 585310 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect 585310 704518 585930 704602
rect 585310 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect 585310 687454 585930 704282
rect 585310 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 585930 687454
rect 585310 687134 585930 687218
rect 585310 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 585930 687134
rect 585310 651454 585930 686898
rect 585310 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 585930 651454
rect 585310 651134 585930 651218
rect 585310 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 585930 651134
rect 585310 615454 585930 650898
rect 585310 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 585930 615454
rect 585310 615134 585930 615218
rect 585310 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 585930 615134
rect 585310 579454 585930 614898
rect 585310 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 585930 579454
rect 585310 579134 585930 579218
rect 585310 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 585930 579134
rect 585310 543454 585930 578898
rect 585310 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 585930 543454
rect 585310 543134 585930 543218
rect 585310 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 585930 543134
rect 585310 507454 585930 542898
rect 585310 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 585930 507454
rect 585310 507134 585930 507218
rect 585310 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 585930 507134
rect 585310 471454 585930 506898
rect 585310 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 585930 471454
rect 585310 471134 585930 471218
rect 585310 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 585930 471134
rect 585310 435454 585930 470898
rect 585310 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 585930 435454
rect 585310 435134 585930 435218
rect 585310 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 585930 435134
rect 585310 399454 585930 434898
rect 585310 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 585930 399454
rect 585310 399134 585930 399218
rect 585310 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 585930 399134
rect 585310 363454 585930 398898
rect 585310 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 585930 363454
rect 585310 363134 585930 363218
rect 585310 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 585930 363134
rect 585310 327454 585930 362898
rect 585310 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 585930 327454
rect 585310 327134 585930 327218
rect 585310 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 585930 327134
rect 585310 291454 585930 326898
rect 585310 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 585930 291454
rect 585310 291134 585930 291218
rect 585310 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 585930 291134
rect 585310 255454 585930 290898
rect 585310 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 585930 255454
rect 585310 255134 585930 255218
rect 585310 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 585930 255134
rect 585310 219454 585930 254898
rect 585310 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 585930 219454
rect 585310 219134 585930 219218
rect 585310 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 585930 219134
rect 585310 183454 585930 218898
rect 585310 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 585930 183454
rect 585310 183134 585930 183218
rect 585310 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 585930 183134
rect 585310 147454 585930 182898
rect 585310 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 585930 147454
rect 585310 147134 585930 147218
rect 585310 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 585930 147134
rect 585310 111454 585930 146898
rect 585310 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 585930 111454
rect 585310 111134 585930 111218
rect 585310 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 585930 111134
rect 585310 75454 585930 110898
rect 585310 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 585930 75454
rect 585310 75134 585930 75218
rect 585310 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 585930 75134
rect 585310 39454 585930 74898
rect 585310 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 585930 39454
rect 585310 39134 585930 39218
rect 585310 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 585930 39134
rect 585310 3454 585930 38898
rect 585310 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 585930 3454
rect 585310 3134 585930 3218
rect 585310 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 585930 3134
rect 585310 -346 585930 2898
rect 585310 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect 585310 -666 585930 -582
rect 585310 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect 585310 -934 585930 -902
rect 586270 669454 586890 705242
rect 586270 669218 586302 669454
rect 586538 669218 586622 669454
rect 586858 669218 586890 669454
rect 586270 669134 586890 669218
rect 586270 668898 586302 669134
rect 586538 668898 586622 669134
rect 586858 668898 586890 669134
rect 586270 633454 586890 668898
rect 586270 633218 586302 633454
rect 586538 633218 586622 633454
rect 586858 633218 586890 633454
rect 586270 633134 586890 633218
rect 586270 632898 586302 633134
rect 586538 632898 586622 633134
rect 586858 632898 586890 633134
rect 586270 597454 586890 632898
rect 586270 597218 586302 597454
rect 586538 597218 586622 597454
rect 586858 597218 586890 597454
rect 586270 597134 586890 597218
rect 586270 596898 586302 597134
rect 586538 596898 586622 597134
rect 586858 596898 586890 597134
rect 586270 561454 586890 596898
rect 586270 561218 586302 561454
rect 586538 561218 586622 561454
rect 586858 561218 586890 561454
rect 586270 561134 586890 561218
rect 586270 560898 586302 561134
rect 586538 560898 586622 561134
rect 586858 560898 586890 561134
rect 586270 525454 586890 560898
rect 586270 525218 586302 525454
rect 586538 525218 586622 525454
rect 586858 525218 586890 525454
rect 586270 525134 586890 525218
rect 586270 524898 586302 525134
rect 586538 524898 586622 525134
rect 586858 524898 586890 525134
rect 586270 489454 586890 524898
rect 586270 489218 586302 489454
rect 586538 489218 586622 489454
rect 586858 489218 586890 489454
rect 586270 489134 586890 489218
rect 586270 488898 586302 489134
rect 586538 488898 586622 489134
rect 586858 488898 586890 489134
rect 586270 453454 586890 488898
rect 586270 453218 586302 453454
rect 586538 453218 586622 453454
rect 586858 453218 586890 453454
rect 586270 453134 586890 453218
rect 586270 452898 586302 453134
rect 586538 452898 586622 453134
rect 586858 452898 586890 453134
rect 586270 417454 586890 452898
rect 586270 417218 586302 417454
rect 586538 417218 586622 417454
rect 586858 417218 586890 417454
rect 586270 417134 586890 417218
rect 586270 416898 586302 417134
rect 586538 416898 586622 417134
rect 586858 416898 586890 417134
rect 586270 381454 586890 416898
rect 586270 381218 586302 381454
rect 586538 381218 586622 381454
rect 586858 381218 586890 381454
rect 586270 381134 586890 381218
rect 586270 380898 586302 381134
rect 586538 380898 586622 381134
rect 586858 380898 586890 381134
rect 586270 345454 586890 380898
rect 586270 345218 586302 345454
rect 586538 345218 586622 345454
rect 586858 345218 586890 345454
rect 586270 345134 586890 345218
rect 586270 344898 586302 345134
rect 586538 344898 586622 345134
rect 586858 344898 586890 345134
rect 586270 309454 586890 344898
rect 586270 309218 586302 309454
rect 586538 309218 586622 309454
rect 586858 309218 586890 309454
rect 586270 309134 586890 309218
rect 586270 308898 586302 309134
rect 586538 308898 586622 309134
rect 586858 308898 586890 309134
rect 586270 273454 586890 308898
rect 586270 273218 586302 273454
rect 586538 273218 586622 273454
rect 586858 273218 586890 273454
rect 586270 273134 586890 273218
rect 586270 272898 586302 273134
rect 586538 272898 586622 273134
rect 586858 272898 586890 273134
rect 586270 237454 586890 272898
rect 586270 237218 586302 237454
rect 586538 237218 586622 237454
rect 586858 237218 586890 237454
rect 586270 237134 586890 237218
rect 586270 236898 586302 237134
rect 586538 236898 586622 237134
rect 586858 236898 586890 237134
rect 586270 201454 586890 236898
rect 586270 201218 586302 201454
rect 586538 201218 586622 201454
rect 586858 201218 586890 201454
rect 586270 201134 586890 201218
rect 586270 200898 586302 201134
rect 586538 200898 586622 201134
rect 586858 200898 586890 201134
rect 586270 165454 586890 200898
rect 586270 165218 586302 165454
rect 586538 165218 586622 165454
rect 586858 165218 586890 165454
rect 586270 165134 586890 165218
rect 586270 164898 586302 165134
rect 586538 164898 586622 165134
rect 586858 164898 586890 165134
rect 586270 129454 586890 164898
rect 586270 129218 586302 129454
rect 586538 129218 586622 129454
rect 586858 129218 586890 129454
rect 586270 129134 586890 129218
rect 586270 128898 586302 129134
rect 586538 128898 586622 129134
rect 586858 128898 586890 129134
rect 586270 93454 586890 128898
rect 586270 93218 586302 93454
rect 586538 93218 586622 93454
rect 586858 93218 586890 93454
rect 586270 93134 586890 93218
rect 586270 92898 586302 93134
rect 586538 92898 586622 93134
rect 586858 92898 586890 93134
rect 586270 57454 586890 92898
rect 586270 57218 586302 57454
rect 586538 57218 586622 57454
rect 586858 57218 586890 57454
rect 586270 57134 586890 57218
rect 586270 56898 586302 57134
rect 586538 56898 586622 57134
rect 586858 56898 586890 57134
rect 586270 21454 586890 56898
rect 586270 21218 586302 21454
rect 586538 21218 586622 21454
rect 586858 21218 586890 21454
rect 586270 21134 586890 21218
rect 586270 20898 586302 21134
rect 586538 20898 586622 21134
rect 586858 20898 586890 21134
rect 586270 -1306 586890 20898
rect 586270 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect 586270 -1626 586890 -1542
rect 586270 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect 586270 -1894 586890 -1862
rect 587230 691174 587850 706202
rect 587230 690938 587262 691174
rect 587498 690938 587582 691174
rect 587818 690938 587850 691174
rect 587230 690854 587850 690938
rect 587230 690618 587262 690854
rect 587498 690618 587582 690854
rect 587818 690618 587850 690854
rect 587230 655174 587850 690618
rect 587230 654938 587262 655174
rect 587498 654938 587582 655174
rect 587818 654938 587850 655174
rect 587230 654854 587850 654938
rect 587230 654618 587262 654854
rect 587498 654618 587582 654854
rect 587818 654618 587850 654854
rect 587230 619174 587850 654618
rect 587230 618938 587262 619174
rect 587498 618938 587582 619174
rect 587818 618938 587850 619174
rect 587230 618854 587850 618938
rect 587230 618618 587262 618854
rect 587498 618618 587582 618854
rect 587818 618618 587850 618854
rect 587230 583174 587850 618618
rect 587230 582938 587262 583174
rect 587498 582938 587582 583174
rect 587818 582938 587850 583174
rect 587230 582854 587850 582938
rect 587230 582618 587262 582854
rect 587498 582618 587582 582854
rect 587818 582618 587850 582854
rect 587230 547174 587850 582618
rect 587230 546938 587262 547174
rect 587498 546938 587582 547174
rect 587818 546938 587850 547174
rect 587230 546854 587850 546938
rect 587230 546618 587262 546854
rect 587498 546618 587582 546854
rect 587818 546618 587850 546854
rect 587230 511174 587850 546618
rect 587230 510938 587262 511174
rect 587498 510938 587582 511174
rect 587818 510938 587850 511174
rect 587230 510854 587850 510938
rect 587230 510618 587262 510854
rect 587498 510618 587582 510854
rect 587818 510618 587850 510854
rect 587230 475174 587850 510618
rect 587230 474938 587262 475174
rect 587498 474938 587582 475174
rect 587818 474938 587850 475174
rect 587230 474854 587850 474938
rect 587230 474618 587262 474854
rect 587498 474618 587582 474854
rect 587818 474618 587850 474854
rect 587230 439174 587850 474618
rect 587230 438938 587262 439174
rect 587498 438938 587582 439174
rect 587818 438938 587850 439174
rect 587230 438854 587850 438938
rect 587230 438618 587262 438854
rect 587498 438618 587582 438854
rect 587818 438618 587850 438854
rect 587230 403174 587850 438618
rect 587230 402938 587262 403174
rect 587498 402938 587582 403174
rect 587818 402938 587850 403174
rect 587230 402854 587850 402938
rect 587230 402618 587262 402854
rect 587498 402618 587582 402854
rect 587818 402618 587850 402854
rect 587230 367174 587850 402618
rect 587230 366938 587262 367174
rect 587498 366938 587582 367174
rect 587818 366938 587850 367174
rect 587230 366854 587850 366938
rect 587230 366618 587262 366854
rect 587498 366618 587582 366854
rect 587818 366618 587850 366854
rect 587230 331174 587850 366618
rect 587230 330938 587262 331174
rect 587498 330938 587582 331174
rect 587818 330938 587850 331174
rect 587230 330854 587850 330938
rect 587230 330618 587262 330854
rect 587498 330618 587582 330854
rect 587818 330618 587850 330854
rect 587230 295174 587850 330618
rect 587230 294938 587262 295174
rect 587498 294938 587582 295174
rect 587818 294938 587850 295174
rect 587230 294854 587850 294938
rect 587230 294618 587262 294854
rect 587498 294618 587582 294854
rect 587818 294618 587850 294854
rect 587230 259174 587850 294618
rect 587230 258938 587262 259174
rect 587498 258938 587582 259174
rect 587818 258938 587850 259174
rect 587230 258854 587850 258938
rect 587230 258618 587262 258854
rect 587498 258618 587582 258854
rect 587818 258618 587850 258854
rect 587230 223174 587850 258618
rect 587230 222938 587262 223174
rect 587498 222938 587582 223174
rect 587818 222938 587850 223174
rect 587230 222854 587850 222938
rect 587230 222618 587262 222854
rect 587498 222618 587582 222854
rect 587818 222618 587850 222854
rect 587230 187174 587850 222618
rect 587230 186938 587262 187174
rect 587498 186938 587582 187174
rect 587818 186938 587850 187174
rect 587230 186854 587850 186938
rect 587230 186618 587262 186854
rect 587498 186618 587582 186854
rect 587818 186618 587850 186854
rect 587230 151174 587850 186618
rect 587230 150938 587262 151174
rect 587498 150938 587582 151174
rect 587818 150938 587850 151174
rect 587230 150854 587850 150938
rect 587230 150618 587262 150854
rect 587498 150618 587582 150854
rect 587818 150618 587850 150854
rect 587230 115174 587850 150618
rect 587230 114938 587262 115174
rect 587498 114938 587582 115174
rect 587818 114938 587850 115174
rect 587230 114854 587850 114938
rect 587230 114618 587262 114854
rect 587498 114618 587582 114854
rect 587818 114618 587850 114854
rect 587230 79174 587850 114618
rect 587230 78938 587262 79174
rect 587498 78938 587582 79174
rect 587818 78938 587850 79174
rect 587230 78854 587850 78938
rect 587230 78618 587262 78854
rect 587498 78618 587582 78854
rect 587818 78618 587850 78854
rect 587230 43174 587850 78618
rect 587230 42938 587262 43174
rect 587498 42938 587582 43174
rect 587818 42938 587850 43174
rect 587230 42854 587850 42938
rect 587230 42618 587262 42854
rect 587498 42618 587582 42854
rect 587818 42618 587850 42854
rect 587230 7174 587850 42618
rect 587230 6938 587262 7174
rect 587498 6938 587582 7174
rect 587818 6938 587850 7174
rect 587230 6854 587850 6938
rect 587230 6618 587262 6854
rect 587498 6618 587582 6854
rect 587818 6618 587850 6854
rect 581514 -2502 581546 -2266
rect 581782 -2502 581866 -2266
rect 582102 -2502 582134 -2266
rect 581514 -2586 582134 -2502
rect 581514 -2822 581546 -2586
rect 581782 -2822 581866 -2586
rect 582102 -2822 582134 -2586
rect 581514 -3814 582134 -2822
rect 587230 -2266 587850 6618
rect 587230 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect 587230 -2586 587850 -2502
rect 587230 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect 587230 -2854 587850 -2822
rect 588190 673174 588810 707162
rect 588190 672938 588222 673174
rect 588458 672938 588542 673174
rect 588778 672938 588810 673174
rect 588190 672854 588810 672938
rect 588190 672618 588222 672854
rect 588458 672618 588542 672854
rect 588778 672618 588810 672854
rect 588190 637174 588810 672618
rect 588190 636938 588222 637174
rect 588458 636938 588542 637174
rect 588778 636938 588810 637174
rect 588190 636854 588810 636938
rect 588190 636618 588222 636854
rect 588458 636618 588542 636854
rect 588778 636618 588810 636854
rect 588190 601174 588810 636618
rect 588190 600938 588222 601174
rect 588458 600938 588542 601174
rect 588778 600938 588810 601174
rect 588190 600854 588810 600938
rect 588190 600618 588222 600854
rect 588458 600618 588542 600854
rect 588778 600618 588810 600854
rect 588190 565174 588810 600618
rect 588190 564938 588222 565174
rect 588458 564938 588542 565174
rect 588778 564938 588810 565174
rect 588190 564854 588810 564938
rect 588190 564618 588222 564854
rect 588458 564618 588542 564854
rect 588778 564618 588810 564854
rect 588190 529174 588810 564618
rect 588190 528938 588222 529174
rect 588458 528938 588542 529174
rect 588778 528938 588810 529174
rect 588190 528854 588810 528938
rect 588190 528618 588222 528854
rect 588458 528618 588542 528854
rect 588778 528618 588810 528854
rect 588190 493174 588810 528618
rect 588190 492938 588222 493174
rect 588458 492938 588542 493174
rect 588778 492938 588810 493174
rect 588190 492854 588810 492938
rect 588190 492618 588222 492854
rect 588458 492618 588542 492854
rect 588778 492618 588810 492854
rect 588190 457174 588810 492618
rect 588190 456938 588222 457174
rect 588458 456938 588542 457174
rect 588778 456938 588810 457174
rect 588190 456854 588810 456938
rect 588190 456618 588222 456854
rect 588458 456618 588542 456854
rect 588778 456618 588810 456854
rect 588190 421174 588810 456618
rect 588190 420938 588222 421174
rect 588458 420938 588542 421174
rect 588778 420938 588810 421174
rect 588190 420854 588810 420938
rect 588190 420618 588222 420854
rect 588458 420618 588542 420854
rect 588778 420618 588810 420854
rect 588190 385174 588810 420618
rect 588190 384938 588222 385174
rect 588458 384938 588542 385174
rect 588778 384938 588810 385174
rect 588190 384854 588810 384938
rect 588190 384618 588222 384854
rect 588458 384618 588542 384854
rect 588778 384618 588810 384854
rect 588190 349174 588810 384618
rect 588190 348938 588222 349174
rect 588458 348938 588542 349174
rect 588778 348938 588810 349174
rect 588190 348854 588810 348938
rect 588190 348618 588222 348854
rect 588458 348618 588542 348854
rect 588778 348618 588810 348854
rect 588190 313174 588810 348618
rect 588190 312938 588222 313174
rect 588458 312938 588542 313174
rect 588778 312938 588810 313174
rect 588190 312854 588810 312938
rect 588190 312618 588222 312854
rect 588458 312618 588542 312854
rect 588778 312618 588810 312854
rect 588190 277174 588810 312618
rect 588190 276938 588222 277174
rect 588458 276938 588542 277174
rect 588778 276938 588810 277174
rect 588190 276854 588810 276938
rect 588190 276618 588222 276854
rect 588458 276618 588542 276854
rect 588778 276618 588810 276854
rect 588190 241174 588810 276618
rect 588190 240938 588222 241174
rect 588458 240938 588542 241174
rect 588778 240938 588810 241174
rect 588190 240854 588810 240938
rect 588190 240618 588222 240854
rect 588458 240618 588542 240854
rect 588778 240618 588810 240854
rect 588190 205174 588810 240618
rect 588190 204938 588222 205174
rect 588458 204938 588542 205174
rect 588778 204938 588810 205174
rect 588190 204854 588810 204938
rect 588190 204618 588222 204854
rect 588458 204618 588542 204854
rect 588778 204618 588810 204854
rect 588190 169174 588810 204618
rect 588190 168938 588222 169174
rect 588458 168938 588542 169174
rect 588778 168938 588810 169174
rect 588190 168854 588810 168938
rect 588190 168618 588222 168854
rect 588458 168618 588542 168854
rect 588778 168618 588810 168854
rect 588190 133174 588810 168618
rect 588190 132938 588222 133174
rect 588458 132938 588542 133174
rect 588778 132938 588810 133174
rect 588190 132854 588810 132938
rect 588190 132618 588222 132854
rect 588458 132618 588542 132854
rect 588778 132618 588810 132854
rect 588190 97174 588810 132618
rect 588190 96938 588222 97174
rect 588458 96938 588542 97174
rect 588778 96938 588810 97174
rect 588190 96854 588810 96938
rect 588190 96618 588222 96854
rect 588458 96618 588542 96854
rect 588778 96618 588810 96854
rect 588190 61174 588810 96618
rect 588190 60938 588222 61174
rect 588458 60938 588542 61174
rect 588778 60938 588810 61174
rect 588190 60854 588810 60938
rect 588190 60618 588222 60854
rect 588458 60618 588542 60854
rect 588778 60618 588810 60854
rect 588190 25174 588810 60618
rect 588190 24938 588222 25174
rect 588458 24938 588542 25174
rect 588778 24938 588810 25174
rect 588190 24854 588810 24938
rect 588190 24618 588222 24854
rect 588458 24618 588542 24854
rect 588778 24618 588810 24854
rect 588190 -3226 588810 24618
rect 588190 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect 588190 -3546 588810 -3462
rect 588190 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect 588190 -3814 588810 -3782
rect 589150 694894 589770 708122
rect 589150 694658 589182 694894
rect 589418 694658 589502 694894
rect 589738 694658 589770 694894
rect 589150 694574 589770 694658
rect 589150 694338 589182 694574
rect 589418 694338 589502 694574
rect 589738 694338 589770 694574
rect 589150 658894 589770 694338
rect 589150 658658 589182 658894
rect 589418 658658 589502 658894
rect 589738 658658 589770 658894
rect 589150 658574 589770 658658
rect 589150 658338 589182 658574
rect 589418 658338 589502 658574
rect 589738 658338 589770 658574
rect 589150 622894 589770 658338
rect 589150 622658 589182 622894
rect 589418 622658 589502 622894
rect 589738 622658 589770 622894
rect 589150 622574 589770 622658
rect 589150 622338 589182 622574
rect 589418 622338 589502 622574
rect 589738 622338 589770 622574
rect 589150 586894 589770 622338
rect 589150 586658 589182 586894
rect 589418 586658 589502 586894
rect 589738 586658 589770 586894
rect 589150 586574 589770 586658
rect 589150 586338 589182 586574
rect 589418 586338 589502 586574
rect 589738 586338 589770 586574
rect 589150 550894 589770 586338
rect 589150 550658 589182 550894
rect 589418 550658 589502 550894
rect 589738 550658 589770 550894
rect 589150 550574 589770 550658
rect 589150 550338 589182 550574
rect 589418 550338 589502 550574
rect 589738 550338 589770 550574
rect 589150 514894 589770 550338
rect 589150 514658 589182 514894
rect 589418 514658 589502 514894
rect 589738 514658 589770 514894
rect 589150 514574 589770 514658
rect 589150 514338 589182 514574
rect 589418 514338 589502 514574
rect 589738 514338 589770 514574
rect 589150 478894 589770 514338
rect 589150 478658 589182 478894
rect 589418 478658 589502 478894
rect 589738 478658 589770 478894
rect 589150 478574 589770 478658
rect 589150 478338 589182 478574
rect 589418 478338 589502 478574
rect 589738 478338 589770 478574
rect 589150 442894 589770 478338
rect 589150 442658 589182 442894
rect 589418 442658 589502 442894
rect 589738 442658 589770 442894
rect 589150 442574 589770 442658
rect 589150 442338 589182 442574
rect 589418 442338 589502 442574
rect 589738 442338 589770 442574
rect 589150 406894 589770 442338
rect 589150 406658 589182 406894
rect 589418 406658 589502 406894
rect 589738 406658 589770 406894
rect 589150 406574 589770 406658
rect 589150 406338 589182 406574
rect 589418 406338 589502 406574
rect 589738 406338 589770 406574
rect 589150 370894 589770 406338
rect 589150 370658 589182 370894
rect 589418 370658 589502 370894
rect 589738 370658 589770 370894
rect 589150 370574 589770 370658
rect 589150 370338 589182 370574
rect 589418 370338 589502 370574
rect 589738 370338 589770 370574
rect 589150 334894 589770 370338
rect 589150 334658 589182 334894
rect 589418 334658 589502 334894
rect 589738 334658 589770 334894
rect 589150 334574 589770 334658
rect 589150 334338 589182 334574
rect 589418 334338 589502 334574
rect 589738 334338 589770 334574
rect 589150 298894 589770 334338
rect 589150 298658 589182 298894
rect 589418 298658 589502 298894
rect 589738 298658 589770 298894
rect 589150 298574 589770 298658
rect 589150 298338 589182 298574
rect 589418 298338 589502 298574
rect 589738 298338 589770 298574
rect 589150 262894 589770 298338
rect 589150 262658 589182 262894
rect 589418 262658 589502 262894
rect 589738 262658 589770 262894
rect 589150 262574 589770 262658
rect 589150 262338 589182 262574
rect 589418 262338 589502 262574
rect 589738 262338 589770 262574
rect 589150 226894 589770 262338
rect 589150 226658 589182 226894
rect 589418 226658 589502 226894
rect 589738 226658 589770 226894
rect 589150 226574 589770 226658
rect 589150 226338 589182 226574
rect 589418 226338 589502 226574
rect 589738 226338 589770 226574
rect 589150 190894 589770 226338
rect 589150 190658 589182 190894
rect 589418 190658 589502 190894
rect 589738 190658 589770 190894
rect 589150 190574 589770 190658
rect 589150 190338 589182 190574
rect 589418 190338 589502 190574
rect 589738 190338 589770 190574
rect 589150 154894 589770 190338
rect 589150 154658 589182 154894
rect 589418 154658 589502 154894
rect 589738 154658 589770 154894
rect 589150 154574 589770 154658
rect 589150 154338 589182 154574
rect 589418 154338 589502 154574
rect 589738 154338 589770 154574
rect 589150 118894 589770 154338
rect 589150 118658 589182 118894
rect 589418 118658 589502 118894
rect 589738 118658 589770 118894
rect 589150 118574 589770 118658
rect 589150 118338 589182 118574
rect 589418 118338 589502 118574
rect 589738 118338 589770 118574
rect 589150 82894 589770 118338
rect 589150 82658 589182 82894
rect 589418 82658 589502 82894
rect 589738 82658 589770 82894
rect 589150 82574 589770 82658
rect 589150 82338 589182 82574
rect 589418 82338 589502 82574
rect 589738 82338 589770 82574
rect 589150 46894 589770 82338
rect 589150 46658 589182 46894
rect 589418 46658 589502 46894
rect 589738 46658 589770 46894
rect 589150 46574 589770 46658
rect 589150 46338 589182 46574
rect 589418 46338 589502 46574
rect 589738 46338 589770 46574
rect 589150 10894 589770 46338
rect 589150 10658 589182 10894
rect 589418 10658 589502 10894
rect 589738 10658 589770 10894
rect 589150 10574 589770 10658
rect 589150 10338 589182 10574
rect 589418 10338 589502 10574
rect 589738 10338 589770 10574
rect 589150 -4186 589770 10338
rect 589150 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect 589150 -4506 589770 -4422
rect 589150 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect 589150 -4774 589770 -4742
rect 590110 676894 590730 709082
rect 590110 676658 590142 676894
rect 590378 676658 590462 676894
rect 590698 676658 590730 676894
rect 590110 676574 590730 676658
rect 590110 676338 590142 676574
rect 590378 676338 590462 676574
rect 590698 676338 590730 676574
rect 590110 640894 590730 676338
rect 590110 640658 590142 640894
rect 590378 640658 590462 640894
rect 590698 640658 590730 640894
rect 590110 640574 590730 640658
rect 590110 640338 590142 640574
rect 590378 640338 590462 640574
rect 590698 640338 590730 640574
rect 590110 604894 590730 640338
rect 590110 604658 590142 604894
rect 590378 604658 590462 604894
rect 590698 604658 590730 604894
rect 590110 604574 590730 604658
rect 590110 604338 590142 604574
rect 590378 604338 590462 604574
rect 590698 604338 590730 604574
rect 590110 568894 590730 604338
rect 590110 568658 590142 568894
rect 590378 568658 590462 568894
rect 590698 568658 590730 568894
rect 590110 568574 590730 568658
rect 590110 568338 590142 568574
rect 590378 568338 590462 568574
rect 590698 568338 590730 568574
rect 590110 532894 590730 568338
rect 590110 532658 590142 532894
rect 590378 532658 590462 532894
rect 590698 532658 590730 532894
rect 590110 532574 590730 532658
rect 590110 532338 590142 532574
rect 590378 532338 590462 532574
rect 590698 532338 590730 532574
rect 590110 496894 590730 532338
rect 590110 496658 590142 496894
rect 590378 496658 590462 496894
rect 590698 496658 590730 496894
rect 590110 496574 590730 496658
rect 590110 496338 590142 496574
rect 590378 496338 590462 496574
rect 590698 496338 590730 496574
rect 590110 460894 590730 496338
rect 590110 460658 590142 460894
rect 590378 460658 590462 460894
rect 590698 460658 590730 460894
rect 590110 460574 590730 460658
rect 590110 460338 590142 460574
rect 590378 460338 590462 460574
rect 590698 460338 590730 460574
rect 590110 424894 590730 460338
rect 590110 424658 590142 424894
rect 590378 424658 590462 424894
rect 590698 424658 590730 424894
rect 590110 424574 590730 424658
rect 590110 424338 590142 424574
rect 590378 424338 590462 424574
rect 590698 424338 590730 424574
rect 590110 388894 590730 424338
rect 590110 388658 590142 388894
rect 590378 388658 590462 388894
rect 590698 388658 590730 388894
rect 590110 388574 590730 388658
rect 590110 388338 590142 388574
rect 590378 388338 590462 388574
rect 590698 388338 590730 388574
rect 590110 352894 590730 388338
rect 590110 352658 590142 352894
rect 590378 352658 590462 352894
rect 590698 352658 590730 352894
rect 590110 352574 590730 352658
rect 590110 352338 590142 352574
rect 590378 352338 590462 352574
rect 590698 352338 590730 352574
rect 590110 316894 590730 352338
rect 590110 316658 590142 316894
rect 590378 316658 590462 316894
rect 590698 316658 590730 316894
rect 590110 316574 590730 316658
rect 590110 316338 590142 316574
rect 590378 316338 590462 316574
rect 590698 316338 590730 316574
rect 590110 280894 590730 316338
rect 590110 280658 590142 280894
rect 590378 280658 590462 280894
rect 590698 280658 590730 280894
rect 590110 280574 590730 280658
rect 590110 280338 590142 280574
rect 590378 280338 590462 280574
rect 590698 280338 590730 280574
rect 590110 244894 590730 280338
rect 590110 244658 590142 244894
rect 590378 244658 590462 244894
rect 590698 244658 590730 244894
rect 590110 244574 590730 244658
rect 590110 244338 590142 244574
rect 590378 244338 590462 244574
rect 590698 244338 590730 244574
rect 590110 208894 590730 244338
rect 590110 208658 590142 208894
rect 590378 208658 590462 208894
rect 590698 208658 590730 208894
rect 590110 208574 590730 208658
rect 590110 208338 590142 208574
rect 590378 208338 590462 208574
rect 590698 208338 590730 208574
rect 590110 172894 590730 208338
rect 590110 172658 590142 172894
rect 590378 172658 590462 172894
rect 590698 172658 590730 172894
rect 590110 172574 590730 172658
rect 590110 172338 590142 172574
rect 590378 172338 590462 172574
rect 590698 172338 590730 172574
rect 590110 136894 590730 172338
rect 590110 136658 590142 136894
rect 590378 136658 590462 136894
rect 590698 136658 590730 136894
rect 590110 136574 590730 136658
rect 590110 136338 590142 136574
rect 590378 136338 590462 136574
rect 590698 136338 590730 136574
rect 590110 100894 590730 136338
rect 590110 100658 590142 100894
rect 590378 100658 590462 100894
rect 590698 100658 590730 100894
rect 590110 100574 590730 100658
rect 590110 100338 590142 100574
rect 590378 100338 590462 100574
rect 590698 100338 590730 100574
rect 590110 64894 590730 100338
rect 590110 64658 590142 64894
rect 590378 64658 590462 64894
rect 590698 64658 590730 64894
rect 590110 64574 590730 64658
rect 590110 64338 590142 64574
rect 590378 64338 590462 64574
rect 590698 64338 590730 64574
rect 590110 28894 590730 64338
rect 590110 28658 590142 28894
rect 590378 28658 590462 28894
rect 590698 28658 590730 28894
rect 590110 28574 590730 28658
rect 590110 28338 590142 28574
rect 590378 28338 590462 28574
rect 590698 28338 590730 28574
rect 590110 -5146 590730 28338
rect 590110 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect 590110 -5466 590730 -5382
rect 590110 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect 590110 -5734 590730 -5702
rect 591070 698614 591690 710042
rect 591070 698378 591102 698614
rect 591338 698378 591422 698614
rect 591658 698378 591690 698614
rect 591070 698294 591690 698378
rect 591070 698058 591102 698294
rect 591338 698058 591422 698294
rect 591658 698058 591690 698294
rect 591070 662614 591690 698058
rect 591070 662378 591102 662614
rect 591338 662378 591422 662614
rect 591658 662378 591690 662614
rect 591070 662294 591690 662378
rect 591070 662058 591102 662294
rect 591338 662058 591422 662294
rect 591658 662058 591690 662294
rect 591070 626614 591690 662058
rect 591070 626378 591102 626614
rect 591338 626378 591422 626614
rect 591658 626378 591690 626614
rect 591070 626294 591690 626378
rect 591070 626058 591102 626294
rect 591338 626058 591422 626294
rect 591658 626058 591690 626294
rect 591070 590614 591690 626058
rect 591070 590378 591102 590614
rect 591338 590378 591422 590614
rect 591658 590378 591690 590614
rect 591070 590294 591690 590378
rect 591070 590058 591102 590294
rect 591338 590058 591422 590294
rect 591658 590058 591690 590294
rect 591070 554614 591690 590058
rect 591070 554378 591102 554614
rect 591338 554378 591422 554614
rect 591658 554378 591690 554614
rect 591070 554294 591690 554378
rect 591070 554058 591102 554294
rect 591338 554058 591422 554294
rect 591658 554058 591690 554294
rect 591070 518614 591690 554058
rect 591070 518378 591102 518614
rect 591338 518378 591422 518614
rect 591658 518378 591690 518614
rect 591070 518294 591690 518378
rect 591070 518058 591102 518294
rect 591338 518058 591422 518294
rect 591658 518058 591690 518294
rect 591070 482614 591690 518058
rect 591070 482378 591102 482614
rect 591338 482378 591422 482614
rect 591658 482378 591690 482614
rect 591070 482294 591690 482378
rect 591070 482058 591102 482294
rect 591338 482058 591422 482294
rect 591658 482058 591690 482294
rect 591070 446614 591690 482058
rect 591070 446378 591102 446614
rect 591338 446378 591422 446614
rect 591658 446378 591690 446614
rect 591070 446294 591690 446378
rect 591070 446058 591102 446294
rect 591338 446058 591422 446294
rect 591658 446058 591690 446294
rect 591070 410614 591690 446058
rect 591070 410378 591102 410614
rect 591338 410378 591422 410614
rect 591658 410378 591690 410614
rect 591070 410294 591690 410378
rect 591070 410058 591102 410294
rect 591338 410058 591422 410294
rect 591658 410058 591690 410294
rect 591070 374614 591690 410058
rect 591070 374378 591102 374614
rect 591338 374378 591422 374614
rect 591658 374378 591690 374614
rect 591070 374294 591690 374378
rect 591070 374058 591102 374294
rect 591338 374058 591422 374294
rect 591658 374058 591690 374294
rect 591070 338614 591690 374058
rect 591070 338378 591102 338614
rect 591338 338378 591422 338614
rect 591658 338378 591690 338614
rect 591070 338294 591690 338378
rect 591070 338058 591102 338294
rect 591338 338058 591422 338294
rect 591658 338058 591690 338294
rect 591070 302614 591690 338058
rect 591070 302378 591102 302614
rect 591338 302378 591422 302614
rect 591658 302378 591690 302614
rect 591070 302294 591690 302378
rect 591070 302058 591102 302294
rect 591338 302058 591422 302294
rect 591658 302058 591690 302294
rect 591070 266614 591690 302058
rect 591070 266378 591102 266614
rect 591338 266378 591422 266614
rect 591658 266378 591690 266614
rect 591070 266294 591690 266378
rect 591070 266058 591102 266294
rect 591338 266058 591422 266294
rect 591658 266058 591690 266294
rect 591070 230614 591690 266058
rect 591070 230378 591102 230614
rect 591338 230378 591422 230614
rect 591658 230378 591690 230614
rect 591070 230294 591690 230378
rect 591070 230058 591102 230294
rect 591338 230058 591422 230294
rect 591658 230058 591690 230294
rect 591070 194614 591690 230058
rect 591070 194378 591102 194614
rect 591338 194378 591422 194614
rect 591658 194378 591690 194614
rect 591070 194294 591690 194378
rect 591070 194058 591102 194294
rect 591338 194058 591422 194294
rect 591658 194058 591690 194294
rect 591070 158614 591690 194058
rect 591070 158378 591102 158614
rect 591338 158378 591422 158614
rect 591658 158378 591690 158614
rect 591070 158294 591690 158378
rect 591070 158058 591102 158294
rect 591338 158058 591422 158294
rect 591658 158058 591690 158294
rect 591070 122614 591690 158058
rect 591070 122378 591102 122614
rect 591338 122378 591422 122614
rect 591658 122378 591690 122614
rect 591070 122294 591690 122378
rect 591070 122058 591102 122294
rect 591338 122058 591422 122294
rect 591658 122058 591690 122294
rect 591070 86614 591690 122058
rect 591070 86378 591102 86614
rect 591338 86378 591422 86614
rect 591658 86378 591690 86614
rect 591070 86294 591690 86378
rect 591070 86058 591102 86294
rect 591338 86058 591422 86294
rect 591658 86058 591690 86294
rect 591070 50614 591690 86058
rect 591070 50378 591102 50614
rect 591338 50378 591422 50614
rect 591658 50378 591690 50614
rect 591070 50294 591690 50378
rect 591070 50058 591102 50294
rect 591338 50058 591422 50294
rect 591658 50058 591690 50294
rect 591070 14614 591690 50058
rect 591070 14378 591102 14614
rect 591338 14378 591422 14614
rect 591658 14378 591690 14614
rect 591070 14294 591690 14378
rect 591070 14058 591102 14294
rect 591338 14058 591422 14294
rect 591658 14058 591690 14294
rect 591070 -6106 591690 14058
rect 591070 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect 591070 -6426 591690 -6342
rect 591070 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect 591070 -6694 591690 -6662
rect 592030 680614 592650 711002
rect 592030 680378 592062 680614
rect 592298 680378 592382 680614
rect 592618 680378 592650 680614
rect 592030 680294 592650 680378
rect 592030 680058 592062 680294
rect 592298 680058 592382 680294
rect 592618 680058 592650 680294
rect 592030 644614 592650 680058
rect 592030 644378 592062 644614
rect 592298 644378 592382 644614
rect 592618 644378 592650 644614
rect 592030 644294 592650 644378
rect 592030 644058 592062 644294
rect 592298 644058 592382 644294
rect 592618 644058 592650 644294
rect 592030 608614 592650 644058
rect 592030 608378 592062 608614
rect 592298 608378 592382 608614
rect 592618 608378 592650 608614
rect 592030 608294 592650 608378
rect 592030 608058 592062 608294
rect 592298 608058 592382 608294
rect 592618 608058 592650 608294
rect 592030 572614 592650 608058
rect 592030 572378 592062 572614
rect 592298 572378 592382 572614
rect 592618 572378 592650 572614
rect 592030 572294 592650 572378
rect 592030 572058 592062 572294
rect 592298 572058 592382 572294
rect 592618 572058 592650 572294
rect 592030 536614 592650 572058
rect 592030 536378 592062 536614
rect 592298 536378 592382 536614
rect 592618 536378 592650 536614
rect 592030 536294 592650 536378
rect 592030 536058 592062 536294
rect 592298 536058 592382 536294
rect 592618 536058 592650 536294
rect 592030 500614 592650 536058
rect 592030 500378 592062 500614
rect 592298 500378 592382 500614
rect 592618 500378 592650 500614
rect 592030 500294 592650 500378
rect 592030 500058 592062 500294
rect 592298 500058 592382 500294
rect 592618 500058 592650 500294
rect 592030 464614 592650 500058
rect 592030 464378 592062 464614
rect 592298 464378 592382 464614
rect 592618 464378 592650 464614
rect 592030 464294 592650 464378
rect 592030 464058 592062 464294
rect 592298 464058 592382 464294
rect 592618 464058 592650 464294
rect 592030 428614 592650 464058
rect 592030 428378 592062 428614
rect 592298 428378 592382 428614
rect 592618 428378 592650 428614
rect 592030 428294 592650 428378
rect 592030 428058 592062 428294
rect 592298 428058 592382 428294
rect 592618 428058 592650 428294
rect 592030 392614 592650 428058
rect 592030 392378 592062 392614
rect 592298 392378 592382 392614
rect 592618 392378 592650 392614
rect 592030 392294 592650 392378
rect 592030 392058 592062 392294
rect 592298 392058 592382 392294
rect 592618 392058 592650 392294
rect 592030 356614 592650 392058
rect 592030 356378 592062 356614
rect 592298 356378 592382 356614
rect 592618 356378 592650 356614
rect 592030 356294 592650 356378
rect 592030 356058 592062 356294
rect 592298 356058 592382 356294
rect 592618 356058 592650 356294
rect 592030 320614 592650 356058
rect 592030 320378 592062 320614
rect 592298 320378 592382 320614
rect 592618 320378 592650 320614
rect 592030 320294 592650 320378
rect 592030 320058 592062 320294
rect 592298 320058 592382 320294
rect 592618 320058 592650 320294
rect 592030 284614 592650 320058
rect 592030 284378 592062 284614
rect 592298 284378 592382 284614
rect 592618 284378 592650 284614
rect 592030 284294 592650 284378
rect 592030 284058 592062 284294
rect 592298 284058 592382 284294
rect 592618 284058 592650 284294
rect 592030 248614 592650 284058
rect 592030 248378 592062 248614
rect 592298 248378 592382 248614
rect 592618 248378 592650 248614
rect 592030 248294 592650 248378
rect 592030 248058 592062 248294
rect 592298 248058 592382 248294
rect 592618 248058 592650 248294
rect 592030 212614 592650 248058
rect 592030 212378 592062 212614
rect 592298 212378 592382 212614
rect 592618 212378 592650 212614
rect 592030 212294 592650 212378
rect 592030 212058 592062 212294
rect 592298 212058 592382 212294
rect 592618 212058 592650 212294
rect 592030 176614 592650 212058
rect 592030 176378 592062 176614
rect 592298 176378 592382 176614
rect 592618 176378 592650 176614
rect 592030 176294 592650 176378
rect 592030 176058 592062 176294
rect 592298 176058 592382 176294
rect 592618 176058 592650 176294
rect 592030 140614 592650 176058
rect 592030 140378 592062 140614
rect 592298 140378 592382 140614
rect 592618 140378 592650 140614
rect 592030 140294 592650 140378
rect 592030 140058 592062 140294
rect 592298 140058 592382 140294
rect 592618 140058 592650 140294
rect 592030 104614 592650 140058
rect 592030 104378 592062 104614
rect 592298 104378 592382 104614
rect 592618 104378 592650 104614
rect 592030 104294 592650 104378
rect 592030 104058 592062 104294
rect 592298 104058 592382 104294
rect 592618 104058 592650 104294
rect 592030 68614 592650 104058
rect 592030 68378 592062 68614
rect 592298 68378 592382 68614
rect 592618 68378 592650 68614
rect 592030 68294 592650 68378
rect 592030 68058 592062 68294
rect 592298 68058 592382 68294
rect 592618 68058 592650 68294
rect 592030 32614 592650 68058
rect 592030 32378 592062 32614
rect 592298 32378 592382 32614
rect 592618 32378 592650 32614
rect 592030 32294 592650 32378
rect 592030 32058 592062 32294
rect 592298 32058 592382 32294
rect 592618 32058 592650 32294
rect 570954 -7302 570986 -7066
rect 571222 -7302 571306 -7066
rect 571542 -7302 571574 -7066
rect 570954 -7386 571574 -7302
rect 570954 -7622 570986 -7386
rect 571222 -7622 571306 -7386
rect 571542 -7622 571574 -7386
rect 570954 -7654 571574 -7622
rect 592030 -7066 592650 32058
rect 592030 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect 592030 -7386 592650 -7302
rect 592030 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect 592030 -7654 592650 -7622
<< via4 >>
rect -8694 711322 -8458 711558
rect -8374 711322 -8138 711558
rect -8694 711002 -8458 711238
rect -8374 711002 -8138 711238
rect -8694 680378 -8458 680614
rect -8374 680378 -8138 680614
rect -8694 680058 -8458 680294
rect -8374 680058 -8138 680294
rect -8694 644378 -8458 644614
rect -8374 644378 -8138 644614
rect -8694 644058 -8458 644294
rect -8374 644058 -8138 644294
rect -8694 608378 -8458 608614
rect -8374 608378 -8138 608614
rect -8694 608058 -8458 608294
rect -8374 608058 -8138 608294
rect -8694 572378 -8458 572614
rect -8374 572378 -8138 572614
rect -8694 572058 -8458 572294
rect -8374 572058 -8138 572294
rect -8694 536378 -8458 536614
rect -8374 536378 -8138 536614
rect -8694 536058 -8458 536294
rect -8374 536058 -8138 536294
rect -8694 500378 -8458 500614
rect -8374 500378 -8138 500614
rect -8694 500058 -8458 500294
rect -8374 500058 -8138 500294
rect -8694 464378 -8458 464614
rect -8374 464378 -8138 464614
rect -8694 464058 -8458 464294
rect -8374 464058 -8138 464294
rect -8694 428378 -8458 428614
rect -8374 428378 -8138 428614
rect -8694 428058 -8458 428294
rect -8374 428058 -8138 428294
rect -8694 392378 -8458 392614
rect -8374 392378 -8138 392614
rect -8694 392058 -8458 392294
rect -8374 392058 -8138 392294
rect -8694 356378 -8458 356614
rect -8374 356378 -8138 356614
rect -8694 356058 -8458 356294
rect -8374 356058 -8138 356294
rect -8694 320378 -8458 320614
rect -8374 320378 -8138 320614
rect -8694 320058 -8458 320294
rect -8374 320058 -8138 320294
rect -8694 284378 -8458 284614
rect -8374 284378 -8138 284614
rect -8694 284058 -8458 284294
rect -8374 284058 -8138 284294
rect -8694 248378 -8458 248614
rect -8374 248378 -8138 248614
rect -8694 248058 -8458 248294
rect -8374 248058 -8138 248294
rect -8694 212378 -8458 212614
rect -8374 212378 -8138 212614
rect -8694 212058 -8458 212294
rect -8374 212058 -8138 212294
rect -8694 176378 -8458 176614
rect -8374 176378 -8138 176614
rect -8694 176058 -8458 176294
rect -8374 176058 -8138 176294
rect -8694 140378 -8458 140614
rect -8374 140378 -8138 140614
rect -8694 140058 -8458 140294
rect -8374 140058 -8138 140294
rect -8694 104378 -8458 104614
rect -8374 104378 -8138 104614
rect -8694 104058 -8458 104294
rect -8374 104058 -8138 104294
rect -8694 68378 -8458 68614
rect -8374 68378 -8138 68614
rect -8694 68058 -8458 68294
rect -8374 68058 -8138 68294
rect -8694 32378 -8458 32614
rect -8374 32378 -8138 32614
rect -8694 32058 -8458 32294
rect -8374 32058 -8138 32294
rect -7734 710362 -7498 710598
rect -7414 710362 -7178 710598
rect -7734 710042 -7498 710278
rect -7414 710042 -7178 710278
rect 12986 710362 13222 710598
rect 13306 710362 13542 710598
rect 12986 710042 13222 710278
rect 13306 710042 13542 710278
rect -7734 698378 -7498 698614
rect -7414 698378 -7178 698614
rect -7734 698058 -7498 698294
rect -7414 698058 -7178 698294
rect -7734 662378 -7498 662614
rect -7414 662378 -7178 662614
rect -7734 662058 -7498 662294
rect -7414 662058 -7178 662294
rect -7734 626378 -7498 626614
rect -7414 626378 -7178 626614
rect -7734 626058 -7498 626294
rect -7414 626058 -7178 626294
rect -7734 590378 -7498 590614
rect -7414 590378 -7178 590614
rect -7734 590058 -7498 590294
rect -7414 590058 -7178 590294
rect -7734 554378 -7498 554614
rect -7414 554378 -7178 554614
rect -7734 554058 -7498 554294
rect -7414 554058 -7178 554294
rect -7734 518378 -7498 518614
rect -7414 518378 -7178 518614
rect -7734 518058 -7498 518294
rect -7414 518058 -7178 518294
rect -7734 482378 -7498 482614
rect -7414 482378 -7178 482614
rect -7734 482058 -7498 482294
rect -7414 482058 -7178 482294
rect -7734 446378 -7498 446614
rect -7414 446378 -7178 446614
rect -7734 446058 -7498 446294
rect -7414 446058 -7178 446294
rect -7734 410378 -7498 410614
rect -7414 410378 -7178 410614
rect -7734 410058 -7498 410294
rect -7414 410058 -7178 410294
rect -7734 374378 -7498 374614
rect -7414 374378 -7178 374614
rect -7734 374058 -7498 374294
rect -7414 374058 -7178 374294
rect -7734 338378 -7498 338614
rect -7414 338378 -7178 338614
rect -7734 338058 -7498 338294
rect -7414 338058 -7178 338294
rect -7734 302378 -7498 302614
rect -7414 302378 -7178 302614
rect -7734 302058 -7498 302294
rect -7414 302058 -7178 302294
rect -7734 266378 -7498 266614
rect -7414 266378 -7178 266614
rect -7734 266058 -7498 266294
rect -7414 266058 -7178 266294
rect -7734 230378 -7498 230614
rect -7414 230378 -7178 230614
rect -7734 230058 -7498 230294
rect -7414 230058 -7178 230294
rect -7734 194378 -7498 194614
rect -7414 194378 -7178 194614
rect -7734 194058 -7498 194294
rect -7414 194058 -7178 194294
rect -7734 158378 -7498 158614
rect -7414 158378 -7178 158614
rect -7734 158058 -7498 158294
rect -7414 158058 -7178 158294
rect -7734 122378 -7498 122614
rect -7414 122378 -7178 122614
rect -7734 122058 -7498 122294
rect -7414 122058 -7178 122294
rect -7734 86378 -7498 86614
rect -7414 86378 -7178 86614
rect -7734 86058 -7498 86294
rect -7414 86058 -7178 86294
rect -7734 50378 -7498 50614
rect -7414 50378 -7178 50614
rect -7734 50058 -7498 50294
rect -7414 50058 -7178 50294
rect -7734 14378 -7498 14614
rect -7414 14378 -7178 14614
rect -7734 14058 -7498 14294
rect -7414 14058 -7178 14294
rect -6774 709402 -6538 709638
rect -6454 709402 -6218 709638
rect -6774 709082 -6538 709318
rect -6454 709082 -6218 709318
rect -6774 676658 -6538 676894
rect -6454 676658 -6218 676894
rect -6774 676338 -6538 676574
rect -6454 676338 -6218 676574
rect -6774 640658 -6538 640894
rect -6454 640658 -6218 640894
rect -6774 640338 -6538 640574
rect -6454 640338 -6218 640574
rect -6774 604658 -6538 604894
rect -6454 604658 -6218 604894
rect -6774 604338 -6538 604574
rect -6454 604338 -6218 604574
rect -6774 568658 -6538 568894
rect -6454 568658 -6218 568894
rect -6774 568338 -6538 568574
rect -6454 568338 -6218 568574
rect -6774 532658 -6538 532894
rect -6454 532658 -6218 532894
rect -6774 532338 -6538 532574
rect -6454 532338 -6218 532574
rect -6774 496658 -6538 496894
rect -6454 496658 -6218 496894
rect -6774 496338 -6538 496574
rect -6454 496338 -6218 496574
rect -6774 460658 -6538 460894
rect -6454 460658 -6218 460894
rect -6774 460338 -6538 460574
rect -6454 460338 -6218 460574
rect -6774 424658 -6538 424894
rect -6454 424658 -6218 424894
rect -6774 424338 -6538 424574
rect -6454 424338 -6218 424574
rect -6774 388658 -6538 388894
rect -6454 388658 -6218 388894
rect -6774 388338 -6538 388574
rect -6454 388338 -6218 388574
rect -6774 352658 -6538 352894
rect -6454 352658 -6218 352894
rect -6774 352338 -6538 352574
rect -6454 352338 -6218 352574
rect -6774 316658 -6538 316894
rect -6454 316658 -6218 316894
rect -6774 316338 -6538 316574
rect -6454 316338 -6218 316574
rect -6774 280658 -6538 280894
rect -6454 280658 -6218 280894
rect -6774 280338 -6538 280574
rect -6454 280338 -6218 280574
rect -6774 244658 -6538 244894
rect -6454 244658 -6218 244894
rect -6774 244338 -6538 244574
rect -6454 244338 -6218 244574
rect -6774 208658 -6538 208894
rect -6454 208658 -6218 208894
rect -6774 208338 -6538 208574
rect -6454 208338 -6218 208574
rect -6774 172658 -6538 172894
rect -6454 172658 -6218 172894
rect -6774 172338 -6538 172574
rect -6454 172338 -6218 172574
rect -6774 136658 -6538 136894
rect -6454 136658 -6218 136894
rect -6774 136338 -6538 136574
rect -6454 136338 -6218 136574
rect -6774 100658 -6538 100894
rect -6454 100658 -6218 100894
rect -6774 100338 -6538 100574
rect -6454 100338 -6218 100574
rect -6774 64658 -6538 64894
rect -6454 64658 -6218 64894
rect -6774 64338 -6538 64574
rect -6454 64338 -6218 64574
rect -6774 28658 -6538 28894
rect -6454 28658 -6218 28894
rect -6774 28338 -6538 28574
rect -6454 28338 -6218 28574
rect -5814 708442 -5578 708678
rect -5494 708442 -5258 708678
rect -5814 708122 -5578 708358
rect -5494 708122 -5258 708358
rect 9266 708442 9502 708678
rect 9586 708442 9822 708678
rect 9266 708122 9502 708358
rect 9586 708122 9822 708358
rect -5814 694658 -5578 694894
rect -5494 694658 -5258 694894
rect -5814 694338 -5578 694574
rect -5494 694338 -5258 694574
rect -5814 658658 -5578 658894
rect -5494 658658 -5258 658894
rect -5814 658338 -5578 658574
rect -5494 658338 -5258 658574
rect -5814 622658 -5578 622894
rect -5494 622658 -5258 622894
rect -5814 622338 -5578 622574
rect -5494 622338 -5258 622574
rect -5814 586658 -5578 586894
rect -5494 586658 -5258 586894
rect -5814 586338 -5578 586574
rect -5494 586338 -5258 586574
rect -5814 550658 -5578 550894
rect -5494 550658 -5258 550894
rect -5814 550338 -5578 550574
rect -5494 550338 -5258 550574
rect -5814 514658 -5578 514894
rect -5494 514658 -5258 514894
rect -5814 514338 -5578 514574
rect -5494 514338 -5258 514574
rect -5814 478658 -5578 478894
rect -5494 478658 -5258 478894
rect -5814 478338 -5578 478574
rect -5494 478338 -5258 478574
rect -5814 442658 -5578 442894
rect -5494 442658 -5258 442894
rect -5814 442338 -5578 442574
rect -5494 442338 -5258 442574
rect -5814 406658 -5578 406894
rect -5494 406658 -5258 406894
rect -5814 406338 -5578 406574
rect -5494 406338 -5258 406574
rect -5814 370658 -5578 370894
rect -5494 370658 -5258 370894
rect -5814 370338 -5578 370574
rect -5494 370338 -5258 370574
rect -5814 334658 -5578 334894
rect -5494 334658 -5258 334894
rect -5814 334338 -5578 334574
rect -5494 334338 -5258 334574
rect -5814 298658 -5578 298894
rect -5494 298658 -5258 298894
rect -5814 298338 -5578 298574
rect -5494 298338 -5258 298574
rect -5814 262658 -5578 262894
rect -5494 262658 -5258 262894
rect -5814 262338 -5578 262574
rect -5494 262338 -5258 262574
rect -5814 226658 -5578 226894
rect -5494 226658 -5258 226894
rect -5814 226338 -5578 226574
rect -5494 226338 -5258 226574
rect -5814 190658 -5578 190894
rect -5494 190658 -5258 190894
rect -5814 190338 -5578 190574
rect -5494 190338 -5258 190574
rect -5814 154658 -5578 154894
rect -5494 154658 -5258 154894
rect -5814 154338 -5578 154574
rect -5494 154338 -5258 154574
rect -5814 118658 -5578 118894
rect -5494 118658 -5258 118894
rect -5814 118338 -5578 118574
rect -5494 118338 -5258 118574
rect -5814 82658 -5578 82894
rect -5494 82658 -5258 82894
rect -5814 82338 -5578 82574
rect -5494 82338 -5258 82574
rect -5814 46658 -5578 46894
rect -5494 46658 -5258 46894
rect -5814 46338 -5578 46574
rect -5494 46338 -5258 46574
rect -5814 10658 -5578 10894
rect -5494 10658 -5258 10894
rect -5814 10338 -5578 10574
rect -5494 10338 -5258 10574
rect -4854 707482 -4618 707718
rect -4534 707482 -4298 707718
rect -4854 707162 -4618 707398
rect -4534 707162 -4298 707398
rect -4854 672938 -4618 673174
rect -4534 672938 -4298 673174
rect -4854 672618 -4618 672854
rect -4534 672618 -4298 672854
rect -4854 636938 -4618 637174
rect -4534 636938 -4298 637174
rect -4854 636618 -4618 636854
rect -4534 636618 -4298 636854
rect -4854 600938 -4618 601174
rect -4534 600938 -4298 601174
rect -4854 600618 -4618 600854
rect -4534 600618 -4298 600854
rect -4854 564938 -4618 565174
rect -4534 564938 -4298 565174
rect -4854 564618 -4618 564854
rect -4534 564618 -4298 564854
rect -4854 528938 -4618 529174
rect -4534 528938 -4298 529174
rect -4854 528618 -4618 528854
rect -4534 528618 -4298 528854
rect -4854 492938 -4618 493174
rect -4534 492938 -4298 493174
rect -4854 492618 -4618 492854
rect -4534 492618 -4298 492854
rect -4854 456938 -4618 457174
rect -4534 456938 -4298 457174
rect -4854 456618 -4618 456854
rect -4534 456618 -4298 456854
rect -4854 420938 -4618 421174
rect -4534 420938 -4298 421174
rect -4854 420618 -4618 420854
rect -4534 420618 -4298 420854
rect -4854 384938 -4618 385174
rect -4534 384938 -4298 385174
rect -4854 384618 -4618 384854
rect -4534 384618 -4298 384854
rect -4854 348938 -4618 349174
rect -4534 348938 -4298 349174
rect -4854 348618 -4618 348854
rect -4534 348618 -4298 348854
rect -4854 312938 -4618 313174
rect -4534 312938 -4298 313174
rect -4854 312618 -4618 312854
rect -4534 312618 -4298 312854
rect -4854 276938 -4618 277174
rect -4534 276938 -4298 277174
rect -4854 276618 -4618 276854
rect -4534 276618 -4298 276854
rect -4854 240938 -4618 241174
rect -4534 240938 -4298 241174
rect -4854 240618 -4618 240854
rect -4534 240618 -4298 240854
rect -4854 204938 -4618 205174
rect -4534 204938 -4298 205174
rect -4854 204618 -4618 204854
rect -4534 204618 -4298 204854
rect -4854 168938 -4618 169174
rect -4534 168938 -4298 169174
rect -4854 168618 -4618 168854
rect -4534 168618 -4298 168854
rect -4854 132938 -4618 133174
rect -4534 132938 -4298 133174
rect -4854 132618 -4618 132854
rect -4534 132618 -4298 132854
rect -4854 96938 -4618 97174
rect -4534 96938 -4298 97174
rect -4854 96618 -4618 96854
rect -4534 96618 -4298 96854
rect -4854 60938 -4618 61174
rect -4534 60938 -4298 61174
rect -4854 60618 -4618 60854
rect -4534 60618 -4298 60854
rect -4854 24938 -4618 25174
rect -4534 24938 -4298 25174
rect -4854 24618 -4618 24854
rect -4534 24618 -4298 24854
rect -3894 706522 -3658 706758
rect -3574 706522 -3338 706758
rect -3894 706202 -3658 706438
rect -3574 706202 -3338 706438
rect 5546 706522 5782 706758
rect 5866 706522 6102 706758
rect 5546 706202 5782 706438
rect 5866 706202 6102 706438
rect -3894 690938 -3658 691174
rect -3574 690938 -3338 691174
rect -3894 690618 -3658 690854
rect -3574 690618 -3338 690854
rect -3894 654938 -3658 655174
rect -3574 654938 -3338 655174
rect -3894 654618 -3658 654854
rect -3574 654618 -3338 654854
rect -3894 618938 -3658 619174
rect -3574 618938 -3338 619174
rect -3894 618618 -3658 618854
rect -3574 618618 -3338 618854
rect -3894 582938 -3658 583174
rect -3574 582938 -3338 583174
rect -3894 582618 -3658 582854
rect -3574 582618 -3338 582854
rect -3894 546938 -3658 547174
rect -3574 546938 -3338 547174
rect -3894 546618 -3658 546854
rect -3574 546618 -3338 546854
rect -3894 510938 -3658 511174
rect -3574 510938 -3338 511174
rect -3894 510618 -3658 510854
rect -3574 510618 -3338 510854
rect -3894 474938 -3658 475174
rect -3574 474938 -3338 475174
rect -3894 474618 -3658 474854
rect -3574 474618 -3338 474854
rect -3894 438938 -3658 439174
rect -3574 438938 -3338 439174
rect -3894 438618 -3658 438854
rect -3574 438618 -3338 438854
rect -3894 402938 -3658 403174
rect -3574 402938 -3338 403174
rect -3894 402618 -3658 402854
rect -3574 402618 -3338 402854
rect -3894 366938 -3658 367174
rect -3574 366938 -3338 367174
rect -3894 366618 -3658 366854
rect -3574 366618 -3338 366854
rect -3894 330938 -3658 331174
rect -3574 330938 -3338 331174
rect -3894 330618 -3658 330854
rect -3574 330618 -3338 330854
rect -3894 294938 -3658 295174
rect -3574 294938 -3338 295174
rect -3894 294618 -3658 294854
rect -3574 294618 -3338 294854
rect -3894 258938 -3658 259174
rect -3574 258938 -3338 259174
rect -3894 258618 -3658 258854
rect -3574 258618 -3338 258854
rect -3894 222938 -3658 223174
rect -3574 222938 -3338 223174
rect -3894 222618 -3658 222854
rect -3574 222618 -3338 222854
rect -3894 186938 -3658 187174
rect -3574 186938 -3338 187174
rect -3894 186618 -3658 186854
rect -3574 186618 -3338 186854
rect -3894 150938 -3658 151174
rect -3574 150938 -3338 151174
rect -3894 150618 -3658 150854
rect -3574 150618 -3338 150854
rect -3894 114938 -3658 115174
rect -3574 114938 -3338 115174
rect -3894 114618 -3658 114854
rect -3574 114618 -3338 114854
rect -3894 78938 -3658 79174
rect -3574 78938 -3338 79174
rect -3894 78618 -3658 78854
rect -3574 78618 -3338 78854
rect -3894 42938 -3658 43174
rect -3574 42938 -3338 43174
rect -3894 42618 -3658 42854
rect -3574 42618 -3338 42854
rect -3894 6938 -3658 7174
rect -3574 6938 -3338 7174
rect -3894 6618 -3658 6854
rect -3574 6618 -3338 6854
rect -2934 705562 -2698 705798
rect -2614 705562 -2378 705798
rect -2934 705242 -2698 705478
rect -2614 705242 -2378 705478
rect -2934 669218 -2698 669454
rect -2614 669218 -2378 669454
rect -2934 668898 -2698 669134
rect -2614 668898 -2378 669134
rect -2934 633218 -2698 633454
rect -2614 633218 -2378 633454
rect -2934 632898 -2698 633134
rect -2614 632898 -2378 633134
rect -2934 597218 -2698 597454
rect -2614 597218 -2378 597454
rect -2934 596898 -2698 597134
rect -2614 596898 -2378 597134
rect -2934 561218 -2698 561454
rect -2614 561218 -2378 561454
rect -2934 560898 -2698 561134
rect -2614 560898 -2378 561134
rect -2934 525218 -2698 525454
rect -2614 525218 -2378 525454
rect -2934 524898 -2698 525134
rect -2614 524898 -2378 525134
rect -2934 489218 -2698 489454
rect -2614 489218 -2378 489454
rect -2934 488898 -2698 489134
rect -2614 488898 -2378 489134
rect -2934 453218 -2698 453454
rect -2614 453218 -2378 453454
rect -2934 452898 -2698 453134
rect -2614 452898 -2378 453134
rect -2934 417218 -2698 417454
rect -2614 417218 -2378 417454
rect -2934 416898 -2698 417134
rect -2614 416898 -2378 417134
rect -2934 381218 -2698 381454
rect -2614 381218 -2378 381454
rect -2934 380898 -2698 381134
rect -2614 380898 -2378 381134
rect -2934 345218 -2698 345454
rect -2614 345218 -2378 345454
rect -2934 344898 -2698 345134
rect -2614 344898 -2378 345134
rect -2934 309218 -2698 309454
rect -2614 309218 -2378 309454
rect -2934 308898 -2698 309134
rect -2614 308898 -2378 309134
rect -2934 273218 -2698 273454
rect -2614 273218 -2378 273454
rect -2934 272898 -2698 273134
rect -2614 272898 -2378 273134
rect -2934 237218 -2698 237454
rect -2614 237218 -2378 237454
rect -2934 236898 -2698 237134
rect -2614 236898 -2378 237134
rect -2934 201218 -2698 201454
rect -2614 201218 -2378 201454
rect -2934 200898 -2698 201134
rect -2614 200898 -2378 201134
rect -2934 165218 -2698 165454
rect -2614 165218 -2378 165454
rect -2934 164898 -2698 165134
rect -2614 164898 -2378 165134
rect -2934 129218 -2698 129454
rect -2614 129218 -2378 129454
rect -2934 128898 -2698 129134
rect -2614 128898 -2378 129134
rect -2934 93218 -2698 93454
rect -2614 93218 -2378 93454
rect -2934 92898 -2698 93134
rect -2614 92898 -2378 93134
rect -2934 57218 -2698 57454
rect -2614 57218 -2378 57454
rect -2934 56898 -2698 57134
rect -2614 56898 -2378 57134
rect -2934 21218 -2698 21454
rect -2614 21218 -2378 21454
rect -2934 20898 -2698 21134
rect -2614 20898 -2378 21134
rect -1974 704602 -1738 704838
rect -1654 704602 -1418 704838
rect -1974 704282 -1738 704518
rect -1654 704282 -1418 704518
rect -1974 687218 -1738 687454
rect -1654 687218 -1418 687454
rect -1974 686898 -1738 687134
rect -1654 686898 -1418 687134
rect -1974 651218 -1738 651454
rect -1654 651218 -1418 651454
rect -1974 650898 -1738 651134
rect -1654 650898 -1418 651134
rect -1974 615218 -1738 615454
rect -1654 615218 -1418 615454
rect -1974 614898 -1738 615134
rect -1654 614898 -1418 615134
rect -1974 579218 -1738 579454
rect -1654 579218 -1418 579454
rect -1974 578898 -1738 579134
rect -1654 578898 -1418 579134
rect -1974 543218 -1738 543454
rect -1654 543218 -1418 543454
rect -1974 542898 -1738 543134
rect -1654 542898 -1418 543134
rect -1974 507218 -1738 507454
rect -1654 507218 -1418 507454
rect -1974 506898 -1738 507134
rect -1654 506898 -1418 507134
rect -1974 471218 -1738 471454
rect -1654 471218 -1418 471454
rect -1974 470898 -1738 471134
rect -1654 470898 -1418 471134
rect -1974 435218 -1738 435454
rect -1654 435218 -1418 435454
rect -1974 434898 -1738 435134
rect -1654 434898 -1418 435134
rect -1974 399218 -1738 399454
rect -1654 399218 -1418 399454
rect -1974 398898 -1738 399134
rect -1654 398898 -1418 399134
rect -1974 363218 -1738 363454
rect -1654 363218 -1418 363454
rect -1974 362898 -1738 363134
rect -1654 362898 -1418 363134
rect -1974 327218 -1738 327454
rect -1654 327218 -1418 327454
rect -1974 326898 -1738 327134
rect -1654 326898 -1418 327134
rect -1974 291218 -1738 291454
rect -1654 291218 -1418 291454
rect -1974 290898 -1738 291134
rect -1654 290898 -1418 291134
rect -1974 255218 -1738 255454
rect -1654 255218 -1418 255454
rect -1974 254898 -1738 255134
rect -1654 254898 -1418 255134
rect -1974 219218 -1738 219454
rect -1654 219218 -1418 219454
rect -1974 218898 -1738 219134
rect -1654 218898 -1418 219134
rect -1974 183218 -1738 183454
rect -1654 183218 -1418 183454
rect -1974 182898 -1738 183134
rect -1654 182898 -1418 183134
rect -1974 147218 -1738 147454
rect -1654 147218 -1418 147454
rect -1974 146898 -1738 147134
rect -1654 146898 -1418 147134
rect -1974 111218 -1738 111454
rect -1654 111218 -1418 111454
rect -1974 110898 -1738 111134
rect -1654 110898 -1418 111134
rect -1974 75218 -1738 75454
rect -1654 75218 -1418 75454
rect -1974 74898 -1738 75134
rect -1654 74898 -1418 75134
rect -1974 39218 -1738 39454
rect -1654 39218 -1418 39454
rect -1974 38898 -1738 39134
rect -1654 38898 -1418 39134
rect -1974 3218 -1738 3454
rect -1654 3218 -1418 3454
rect -1974 2898 -1738 3134
rect -1654 2898 -1418 3134
rect -1974 -582 -1738 -346
rect -1654 -582 -1418 -346
rect -1974 -902 -1738 -666
rect -1654 -902 -1418 -666
rect 1826 704602 2062 704838
rect 2146 704602 2382 704838
rect 1826 704282 2062 704518
rect 2146 704282 2382 704518
rect 1826 687218 2062 687454
rect 2146 687218 2382 687454
rect 1826 686898 2062 687134
rect 2146 686898 2382 687134
rect 1826 651218 2062 651454
rect 2146 651218 2382 651454
rect 1826 650898 2062 651134
rect 2146 650898 2382 651134
rect 1826 615218 2062 615454
rect 2146 615218 2382 615454
rect 1826 614898 2062 615134
rect 2146 614898 2382 615134
rect 1826 579218 2062 579454
rect 2146 579218 2382 579454
rect 1826 578898 2062 579134
rect 2146 578898 2382 579134
rect 1826 543218 2062 543454
rect 2146 543218 2382 543454
rect 1826 542898 2062 543134
rect 2146 542898 2382 543134
rect 1826 507218 2062 507454
rect 2146 507218 2382 507454
rect 1826 506898 2062 507134
rect 2146 506898 2382 507134
rect 1826 471218 2062 471454
rect 2146 471218 2382 471454
rect 1826 470898 2062 471134
rect 2146 470898 2382 471134
rect 1826 435218 2062 435454
rect 2146 435218 2382 435454
rect 1826 434898 2062 435134
rect 2146 434898 2382 435134
rect 1826 399218 2062 399454
rect 2146 399218 2382 399454
rect 1826 398898 2062 399134
rect 2146 398898 2382 399134
rect 1826 363218 2062 363454
rect 2146 363218 2382 363454
rect 1826 362898 2062 363134
rect 2146 362898 2382 363134
rect 1826 327218 2062 327454
rect 2146 327218 2382 327454
rect 1826 326898 2062 327134
rect 2146 326898 2382 327134
rect 1826 291218 2062 291454
rect 2146 291218 2382 291454
rect 1826 290898 2062 291134
rect 2146 290898 2382 291134
rect 1826 255218 2062 255454
rect 2146 255218 2382 255454
rect 1826 254898 2062 255134
rect 2146 254898 2382 255134
rect 1826 219218 2062 219454
rect 2146 219218 2382 219454
rect 1826 218898 2062 219134
rect 2146 218898 2382 219134
rect 1826 183218 2062 183454
rect 2146 183218 2382 183454
rect 1826 182898 2062 183134
rect 2146 182898 2382 183134
rect 1826 147218 2062 147454
rect 2146 147218 2382 147454
rect 1826 146898 2062 147134
rect 2146 146898 2382 147134
rect 1826 111218 2062 111454
rect 2146 111218 2382 111454
rect 1826 110898 2062 111134
rect 2146 110898 2382 111134
rect 1826 75218 2062 75454
rect 2146 75218 2382 75454
rect 1826 74898 2062 75134
rect 2146 74898 2382 75134
rect 1826 39218 2062 39454
rect 2146 39218 2382 39454
rect 1826 38898 2062 39134
rect 2146 38898 2382 39134
rect 1826 3218 2062 3454
rect 2146 3218 2382 3454
rect 1826 2898 2062 3134
rect 2146 2898 2382 3134
rect 1826 -582 2062 -346
rect 2146 -582 2382 -346
rect 1826 -902 2062 -666
rect 2146 -902 2382 -666
rect -2934 -1542 -2698 -1306
rect -2614 -1542 -2378 -1306
rect -2934 -1862 -2698 -1626
rect -2614 -1862 -2378 -1626
rect 5546 690938 5782 691174
rect 5866 690938 6102 691174
rect 5546 690618 5782 690854
rect 5866 690618 6102 690854
rect 5546 654938 5782 655174
rect 5866 654938 6102 655174
rect 5546 654618 5782 654854
rect 5866 654618 6102 654854
rect 5546 618938 5782 619174
rect 5866 618938 6102 619174
rect 5546 618618 5782 618854
rect 5866 618618 6102 618854
rect 5546 582938 5782 583174
rect 5866 582938 6102 583174
rect 5546 582618 5782 582854
rect 5866 582618 6102 582854
rect 5546 546938 5782 547174
rect 5866 546938 6102 547174
rect 5546 546618 5782 546854
rect 5866 546618 6102 546854
rect 5546 510938 5782 511174
rect 5866 510938 6102 511174
rect 5546 510618 5782 510854
rect 5866 510618 6102 510854
rect 5546 474938 5782 475174
rect 5866 474938 6102 475174
rect 5546 474618 5782 474854
rect 5866 474618 6102 474854
rect 5546 438938 5782 439174
rect 5866 438938 6102 439174
rect 5546 438618 5782 438854
rect 5866 438618 6102 438854
rect 5546 402938 5782 403174
rect 5866 402938 6102 403174
rect 5546 402618 5782 402854
rect 5866 402618 6102 402854
rect 5546 366938 5782 367174
rect 5866 366938 6102 367174
rect 5546 366618 5782 366854
rect 5866 366618 6102 366854
rect 5546 330938 5782 331174
rect 5866 330938 6102 331174
rect 5546 330618 5782 330854
rect 5866 330618 6102 330854
rect 5546 294938 5782 295174
rect 5866 294938 6102 295174
rect 5546 294618 5782 294854
rect 5866 294618 6102 294854
rect 5546 258938 5782 259174
rect 5866 258938 6102 259174
rect 5546 258618 5782 258854
rect 5866 258618 6102 258854
rect 5546 222938 5782 223174
rect 5866 222938 6102 223174
rect 5546 222618 5782 222854
rect 5866 222618 6102 222854
rect 5546 186938 5782 187174
rect 5866 186938 6102 187174
rect 5546 186618 5782 186854
rect 5866 186618 6102 186854
rect 5546 150938 5782 151174
rect 5866 150938 6102 151174
rect 5546 150618 5782 150854
rect 5866 150618 6102 150854
rect 5546 114938 5782 115174
rect 5866 114938 6102 115174
rect 5546 114618 5782 114854
rect 5866 114618 6102 114854
rect 5546 78938 5782 79174
rect 5866 78938 6102 79174
rect 5546 78618 5782 78854
rect 5866 78618 6102 78854
rect 5546 42938 5782 43174
rect 5866 42938 6102 43174
rect 5546 42618 5782 42854
rect 5866 42618 6102 42854
rect 5546 6938 5782 7174
rect 5866 6938 6102 7174
rect 5546 6618 5782 6854
rect 5866 6618 6102 6854
rect -3894 -2502 -3658 -2266
rect -3574 -2502 -3338 -2266
rect -3894 -2822 -3658 -2586
rect -3574 -2822 -3338 -2586
rect 5546 -2502 5782 -2266
rect 5866 -2502 6102 -2266
rect 5546 -2822 5782 -2586
rect 5866 -2822 6102 -2586
rect -4854 -3462 -4618 -3226
rect -4534 -3462 -4298 -3226
rect -4854 -3782 -4618 -3546
rect -4534 -3782 -4298 -3546
rect 9266 694658 9502 694894
rect 9586 694658 9822 694894
rect 9266 694338 9502 694574
rect 9586 694338 9822 694574
rect 9266 658658 9502 658894
rect 9586 658658 9822 658894
rect 9266 658338 9502 658574
rect 9586 658338 9822 658574
rect 9266 622658 9502 622894
rect 9586 622658 9822 622894
rect 9266 622338 9502 622574
rect 9586 622338 9822 622574
rect 9266 586658 9502 586894
rect 9586 586658 9822 586894
rect 9266 586338 9502 586574
rect 9586 586338 9822 586574
rect 9266 550658 9502 550894
rect 9586 550658 9822 550894
rect 9266 550338 9502 550574
rect 9586 550338 9822 550574
rect 9266 514658 9502 514894
rect 9586 514658 9822 514894
rect 9266 514338 9502 514574
rect 9586 514338 9822 514574
rect 9266 478658 9502 478894
rect 9586 478658 9822 478894
rect 9266 478338 9502 478574
rect 9586 478338 9822 478574
rect 9266 442658 9502 442894
rect 9586 442658 9822 442894
rect 9266 442338 9502 442574
rect 9586 442338 9822 442574
rect 9266 406658 9502 406894
rect 9586 406658 9822 406894
rect 9266 406338 9502 406574
rect 9586 406338 9822 406574
rect 9266 370658 9502 370894
rect 9586 370658 9822 370894
rect 9266 370338 9502 370574
rect 9586 370338 9822 370574
rect 9266 334658 9502 334894
rect 9586 334658 9822 334894
rect 9266 334338 9502 334574
rect 9586 334338 9822 334574
rect 9266 298658 9502 298894
rect 9586 298658 9822 298894
rect 9266 298338 9502 298574
rect 9586 298338 9822 298574
rect 9266 262658 9502 262894
rect 9586 262658 9822 262894
rect 9266 262338 9502 262574
rect 9586 262338 9822 262574
rect 9266 226658 9502 226894
rect 9586 226658 9822 226894
rect 9266 226338 9502 226574
rect 9586 226338 9822 226574
rect 9266 190658 9502 190894
rect 9586 190658 9822 190894
rect 9266 190338 9502 190574
rect 9586 190338 9822 190574
rect 9266 154658 9502 154894
rect 9586 154658 9822 154894
rect 9266 154338 9502 154574
rect 9586 154338 9822 154574
rect 9266 118658 9502 118894
rect 9586 118658 9822 118894
rect 9266 118338 9502 118574
rect 9586 118338 9822 118574
rect 9266 82658 9502 82894
rect 9586 82658 9822 82894
rect 9266 82338 9502 82574
rect 9586 82338 9822 82574
rect 9266 46658 9502 46894
rect 9586 46658 9822 46894
rect 9266 46338 9502 46574
rect 9586 46338 9822 46574
rect 9266 10658 9502 10894
rect 9586 10658 9822 10894
rect 9266 10338 9502 10574
rect 9586 10338 9822 10574
rect -5814 -4422 -5578 -4186
rect -5494 -4422 -5258 -4186
rect -5814 -4742 -5578 -4506
rect -5494 -4742 -5258 -4506
rect 9266 -4422 9502 -4186
rect 9586 -4422 9822 -4186
rect 9266 -4742 9502 -4506
rect 9586 -4742 9822 -4506
rect -6774 -5382 -6538 -5146
rect -6454 -5382 -6218 -5146
rect -6774 -5702 -6538 -5466
rect -6454 -5702 -6218 -5466
rect 30986 711322 31222 711558
rect 31306 711322 31542 711558
rect 30986 711002 31222 711238
rect 31306 711002 31542 711238
rect 27266 709402 27502 709638
rect 27586 709402 27822 709638
rect 27266 709082 27502 709318
rect 27586 709082 27822 709318
rect 23546 707482 23782 707718
rect 23866 707482 24102 707718
rect 23546 707162 23782 707398
rect 23866 707162 24102 707398
rect 12986 698378 13222 698614
rect 13306 698378 13542 698614
rect 12986 698058 13222 698294
rect 13306 698058 13542 698294
rect 12986 662378 13222 662614
rect 13306 662378 13542 662614
rect 12986 662058 13222 662294
rect 13306 662058 13542 662294
rect 12986 626378 13222 626614
rect 13306 626378 13542 626614
rect 12986 626058 13222 626294
rect 13306 626058 13542 626294
rect 12986 590378 13222 590614
rect 13306 590378 13542 590614
rect 12986 590058 13222 590294
rect 13306 590058 13542 590294
rect 12986 554378 13222 554614
rect 13306 554378 13542 554614
rect 12986 554058 13222 554294
rect 13306 554058 13542 554294
rect 12986 518378 13222 518614
rect 13306 518378 13542 518614
rect 12986 518058 13222 518294
rect 13306 518058 13542 518294
rect 12986 482378 13222 482614
rect 13306 482378 13542 482614
rect 12986 482058 13222 482294
rect 13306 482058 13542 482294
rect 12986 446378 13222 446614
rect 13306 446378 13542 446614
rect 12986 446058 13222 446294
rect 13306 446058 13542 446294
rect 12986 410378 13222 410614
rect 13306 410378 13542 410614
rect 12986 410058 13222 410294
rect 13306 410058 13542 410294
rect 12986 374378 13222 374614
rect 13306 374378 13542 374614
rect 12986 374058 13222 374294
rect 13306 374058 13542 374294
rect 12986 338378 13222 338614
rect 13306 338378 13542 338614
rect 12986 338058 13222 338294
rect 13306 338058 13542 338294
rect 12986 302378 13222 302614
rect 13306 302378 13542 302614
rect 12986 302058 13222 302294
rect 13306 302058 13542 302294
rect 12986 266378 13222 266614
rect 13306 266378 13542 266614
rect 12986 266058 13222 266294
rect 13306 266058 13542 266294
rect 12986 230378 13222 230614
rect 13306 230378 13542 230614
rect 12986 230058 13222 230294
rect 13306 230058 13542 230294
rect 12986 194378 13222 194614
rect 13306 194378 13542 194614
rect 12986 194058 13222 194294
rect 13306 194058 13542 194294
rect 12986 158378 13222 158614
rect 13306 158378 13542 158614
rect 12986 158058 13222 158294
rect 13306 158058 13542 158294
rect 12986 122378 13222 122614
rect 13306 122378 13542 122614
rect 12986 122058 13222 122294
rect 13306 122058 13542 122294
rect 12986 86378 13222 86614
rect 13306 86378 13542 86614
rect 12986 86058 13222 86294
rect 13306 86058 13542 86294
rect 12986 50378 13222 50614
rect 13306 50378 13542 50614
rect 12986 50058 13222 50294
rect 13306 50058 13542 50294
rect 12986 14378 13222 14614
rect 13306 14378 13542 14614
rect 12986 14058 13222 14294
rect 13306 14058 13542 14294
rect -7734 -6342 -7498 -6106
rect -7414 -6342 -7178 -6106
rect -7734 -6662 -7498 -6426
rect -7414 -6662 -7178 -6426
rect 19826 705562 20062 705798
rect 20146 705562 20382 705798
rect 19826 705242 20062 705478
rect 20146 705242 20382 705478
rect 19826 669218 20062 669454
rect 20146 669218 20382 669454
rect 19826 668898 20062 669134
rect 20146 668898 20382 669134
rect 19826 633218 20062 633454
rect 20146 633218 20382 633454
rect 19826 632898 20062 633134
rect 20146 632898 20382 633134
rect 19826 597218 20062 597454
rect 20146 597218 20382 597454
rect 19826 596898 20062 597134
rect 20146 596898 20382 597134
rect 19826 561218 20062 561454
rect 20146 561218 20382 561454
rect 19826 560898 20062 561134
rect 20146 560898 20382 561134
rect 19826 525218 20062 525454
rect 20146 525218 20382 525454
rect 19826 524898 20062 525134
rect 20146 524898 20382 525134
rect 19826 489218 20062 489454
rect 20146 489218 20382 489454
rect 19826 488898 20062 489134
rect 20146 488898 20382 489134
rect 19826 453218 20062 453454
rect 20146 453218 20382 453454
rect 19826 452898 20062 453134
rect 20146 452898 20382 453134
rect 19826 417218 20062 417454
rect 20146 417218 20382 417454
rect 19826 416898 20062 417134
rect 20146 416898 20382 417134
rect 19826 381218 20062 381454
rect 20146 381218 20382 381454
rect 19826 380898 20062 381134
rect 20146 380898 20382 381134
rect 19826 345218 20062 345454
rect 20146 345218 20382 345454
rect 19826 344898 20062 345134
rect 20146 344898 20382 345134
rect 19826 309218 20062 309454
rect 20146 309218 20382 309454
rect 19826 308898 20062 309134
rect 20146 308898 20382 309134
rect 19826 273218 20062 273454
rect 20146 273218 20382 273454
rect 19826 272898 20062 273134
rect 20146 272898 20382 273134
rect 19826 237218 20062 237454
rect 20146 237218 20382 237454
rect 19826 236898 20062 237134
rect 20146 236898 20382 237134
rect 19826 201218 20062 201454
rect 20146 201218 20382 201454
rect 19826 200898 20062 201134
rect 20146 200898 20382 201134
rect 19826 165218 20062 165454
rect 20146 165218 20382 165454
rect 19826 164898 20062 165134
rect 20146 164898 20382 165134
rect 19826 129218 20062 129454
rect 20146 129218 20382 129454
rect 19826 128898 20062 129134
rect 20146 128898 20382 129134
rect 19826 93218 20062 93454
rect 20146 93218 20382 93454
rect 19826 92898 20062 93134
rect 20146 92898 20382 93134
rect 19826 57218 20062 57454
rect 20146 57218 20382 57454
rect 19826 56898 20062 57134
rect 20146 56898 20382 57134
rect 19826 21218 20062 21454
rect 20146 21218 20382 21454
rect 19826 20898 20062 21134
rect 20146 20898 20382 21134
rect 19826 -1542 20062 -1306
rect 20146 -1542 20382 -1306
rect 19826 -1862 20062 -1626
rect 20146 -1862 20382 -1626
rect 23546 672938 23782 673174
rect 23866 672938 24102 673174
rect 23546 672618 23782 672854
rect 23866 672618 24102 672854
rect 23546 636938 23782 637174
rect 23866 636938 24102 637174
rect 23546 636618 23782 636854
rect 23866 636618 24102 636854
rect 23546 600938 23782 601174
rect 23866 600938 24102 601174
rect 23546 600618 23782 600854
rect 23866 600618 24102 600854
rect 23546 564938 23782 565174
rect 23866 564938 24102 565174
rect 23546 564618 23782 564854
rect 23866 564618 24102 564854
rect 23546 528938 23782 529174
rect 23866 528938 24102 529174
rect 23546 528618 23782 528854
rect 23866 528618 24102 528854
rect 23546 492938 23782 493174
rect 23866 492938 24102 493174
rect 23546 492618 23782 492854
rect 23866 492618 24102 492854
rect 23546 456938 23782 457174
rect 23866 456938 24102 457174
rect 23546 456618 23782 456854
rect 23866 456618 24102 456854
rect 23546 420938 23782 421174
rect 23866 420938 24102 421174
rect 23546 420618 23782 420854
rect 23866 420618 24102 420854
rect 23546 384938 23782 385174
rect 23866 384938 24102 385174
rect 23546 384618 23782 384854
rect 23866 384618 24102 384854
rect 23546 348938 23782 349174
rect 23866 348938 24102 349174
rect 23546 348618 23782 348854
rect 23866 348618 24102 348854
rect 23546 312938 23782 313174
rect 23866 312938 24102 313174
rect 23546 312618 23782 312854
rect 23866 312618 24102 312854
rect 23546 276938 23782 277174
rect 23866 276938 24102 277174
rect 23546 276618 23782 276854
rect 23866 276618 24102 276854
rect 23546 240938 23782 241174
rect 23866 240938 24102 241174
rect 23546 240618 23782 240854
rect 23866 240618 24102 240854
rect 23546 204938 23782 205174
rect 23866 204938 24102 205174
rect 23546 204618 23782 204854
rect 23866 204618 24102 204854
rect 23546 168938 23782 169174
rect 23866 168938 24102 169174
rect 23546 168618 23782 168854
rect 23866 168618 24102 168854
rect 23546 132938 23782 133174
rect 23866 132938 24102 133174
rect 23546 132618 23782 132854
rect 23866 132618 24102 132854
rect 23546 96938 23782 97174
rect 23866 96938 24102 97174
rect 23546 96618 23782 96854
rect 23866 96618 24102 96854
rect 23546 60938 23782 61174
rect 23866 60938 24102 61174
rect 23546 60618 23782 60854
rect 23866 60618 24102 60854
rect 23546 24938 23782 25174
rect 23866 24938 24102 25174
rect 23546 24618 23782 24854
rect 23866 24618 24102 24854
rect 23546 -3462 23782 -3226
rect 23866 -3462 24102 -3226
rect 23546 -3782 23782 -3546
rect 23866 -3782 24102 -3546
rect 27266 676658 27502 676894
rect 27586 676658 27822 676894
rect 27266 676338 27502 676574
rect 27586 676338 27822 676574
rect 27266 640658 27502 640894
rect 27586 640658 27822 640894
rect 27266 640338 27502 640574
rect 27586 640338 27822 640574
rect 27266 604658 27502 604894
rect 27586 604658 27822 604894
rect 27266 604338 27502 604574
rect 27586 604338 27822 604574
rect 27266 568658 27502 568894
rect 27586 568658 27822 568894
rect 27266 568338 27502 568574
rect 27586 568338 27822 568574
rect 27266 532658 27502 532894
rect 27586 532658 27822 532894
rect 27266 532338 27502 532574
rect 27586 532338 27822 532574
rect 27266 496658 27502 496894
rect 27586 496658 27822 496894
rect 27266 496338 27502 496574
rect 27586 496338 27822 496574
rect 27266 460658 27502 460894
rect 27586 460658 27822 460894
rect 27266 460338 27502 460574
rect 27586 460338 27822 460574
rect 27266 424658 27502 424894
rect 27586 424658 27822 424894
rect 27266 424338 27502 424574
rect 27586 424338 27822 424574
rect 27266 388658 27502 388894
rect 27586 388658 27822 388894
rect 27266 388338 27502 388574
rect 27586 388338 27822 388574
rect 27266 352658 27502 352894
rect 27586 352658 27822 352894
rect 27266 352338 27502 352574
rect 27586 352338 27822 352574
rect 27266 316658 27502 316894
rect 27586 316658 27822 316894
rect 27266 316338 27502 316574
rect 27586 316338 27822 316574
rect 27266 280658 27502 280894
rect 27586 280658 27822 280894
rect 27266 280338 27502 280574
rect 27586 280338 27822 280574
rect 27266 244658 27502 244894
rect 27586 244658 27822 244894
rect 27266 244338 27502 244574
rect 27586 244338 27822 244574
rect 27266 208658 27502 208894
rect 27586 208658 27822 208894
rect 27266 208338 27502 208574
rect 27586 208338 27822 208574
rect 27266 172658 27502 172894
rect 27586 172658 27822 172894
rect 27266 172338 27502 172574
rect 27586 172338 27822 172574
rect 27266 136658 27502 136894
rect 27586 136658 27822 136894
rect 27266 136338 27502 136574
rect 27586 136338 27822 136574
rect 27266 100658 27502 100894
rect 27586 100658 27822 100894
rect 27266 100338 27502 100574
rect 27586 100338 27822 100574
rect 27266 64658 27502 64894
rect 27586 64658 27822 64894
rect 27266 64338 27502 64574
rect 27586 64338 27822 64574
rect 27266 28658 27502 28894
rect 27586 28658 27822 28894
rect 27266 28338 27502 28574
rect 27586 28338 27822 28574
rect 27266 -5382 27502 -5146
rect 27586 -5382 27822 -5146
rect 27266 -5702 27502 -5466
rect 27586 -5702 27822 -5466
rect 48986 710362 49222 710598
rect 49306 710362 49542 710598
rect 48986 710042 49222 710278
rect 49306 710042 49542 710278
rect 45266 708442 45502 708678
rect 45586 708442 45822 708678
rect 45266 708122 45502 708358
rect 45586 708122 45822 708358
rect 41546 706522 41782 706758
rect 41866 706522 42102 706758
rect 41546 706202 41782 706438
rect 41866 706202 42102 706438
rect 30986 680378 31222 680614
rect 31306 680378 31542 680614
rect 30986 680058 31222 680294
rect 31306 680058 31542 680294
rect 30986 644378 31222 644614
rect 31306 644378 31542 644614
rect 30986 644058 31222 644294
rect 31306 644058 31542 644294
rect 30986 608378 31222 608614
rect 31306 608378 31542 608614
rect 30986 608058 31222 608294
rect 31306 608058 31542 608294
rect 30986 572378 31222 572614
rect 31306 572378 31542 572614
rect 30986 572058 31222 572294
rect 31306 572058 31542 572294
rect 30986 536378 31222 536614
rect 31306 536378 31542 536614
rect 30986 536058 31222 536294
rect 31306 536058 31542 536294
rect 30986 500378 31222 500614
rect 31306 500378 31542 500614
rect 30986 500058 31222 500294
rect 31306 500058 31542 500294
rect 30986 464378 31222 464614
rect 31306 464378 31542 464614
rect 30986 464058 31222 464294
rect 31306 464058 31542 464294
rect 30986 428378 31222 428614
rect 31306 428378 31542 428614
rect 30986 428058 31222 428294
rect 31306 428058 31542 428294
rect 30986 392378 31222 392614
rect 31306 392378 31542 392614
rect 30986 392058 31222 392294
rect 31306 392058 31542 392294
rect 30986 356378 31222 356614
rect 31306 356378 31542 356614
rect 30986 356058 31222 356294
rect 31306 356058 31542 356294
rect 30986 320378 31222 320614
rect 31306 320378 31542 320614
rect 30986 320058 31222 320294
rect 31306 320058 31542 320294
rect 30986 284378 31222 284614
rect 31306 284378 31542 284614
rect 30986 284058 31222 284294
rect 31306 284058 31542 284294
rect 30986 248378 31222 248614
rect 31306 248378 31542 248614
rect 30986 248058 31222 248294
rect 31306 248058 31542 248294
rect 30986 212378 31222 212614
rect 31306 212378 31542 212614
rect 30986 212058 31222 212294
rect 31306 212058 31542 212294
rect 30986 176378 31222 176614
rect 31306 176378 31542 176614
rect 30986 176058 31222 176294
rect 31306 176058 31542 176294
rect 30986 140378 31222 140614
rect 31306 140378 31542 140614
rect 30986 140058 31222 140294
rect 31306 140058 31542 140294
rect 30986 104378 31222 104614
rect 31306 104378 31542 104614
rect 30986 104058 31222 104294
rect 31306 104058 31542 104294
rect 30986 68378 31222 68614
rect 31306 68378 31542 68614
rect 30986 68058 31222 68294
rect 31306 68058 31542 68294
rect 30986 32378 31222 32614
rect 31306 32378 31542 32614
rect 30986 32058 31222 32294
rect 31306 32058 31542 32294
rect 12986 -6342 13222 -6106
rect 13306 -6342 13542 -6106
rect 12986 -6662 13222 -6426
rect 13306 -6662 13542 -6426
rect -8694 -7302 -8458 -7066
rect -8374 -7302 -8138 -7066
rect -8694 -7622 -8458 -7386
rect -8374 -7622 -8138 -7386
rect 37826 704602 38062 704838
rect 38146 704602 38382 704838
rect 37826 704282 38062 704518
rect 38146 704282 38382 704518
rect 37826 687218 38062 687454
rect 38146 687218 38382 687454
rect 37826 686898 38062 687134
rect 38146 686898 38382 687134
rect 37826 651218 38062 651454
rect 38146 651218 38382 651454
rect 37826 650898 38062 651134
rect 38146 650898 38382 651134
rect 37826 615218 38062 615454
rect 38146 615218 38382 615454
rect 37826 614898 38062 615134
rect 38146 614898 38382 615134
rect 37826 579218 38062 579454
rect 38146 579218 38382 579454
rect 37826 578898 38062 579134
rect 38146 578898 38382 579134
rect 37826 543218 38062 543454
rect 38146 543218 38382 543454
rect 37826 542898 38062 543134
rect 38146 542898 38382 543134
rect 37826 507218 38062 507454
rect 38146 507218 38382 507454
rect 37826 506898 38062 507134
rect 38146 506898 38382 507134
rect 37826 471218 38062 471454
rect 38146 471218 38382 471454
rect 37826 470898 38062 471134
rect 38146 470898 38382 471134
rect 37826 435218 38062 435454
rect 38146 435218 38382 435454
rect 37826 434898 38062 435134
rect 38146 434898 38382 435134
rect 37826 399218 38062 399454
rect 38146 399218 38382 399454
rect 37826 398898 38062 399134
rect 38146 398898 38382 399134
rect 37826 363218 38062 363454
rect 38146 363218 38382 363454
rect 37826 362898 38062 363134
rect 38146 362898 38382 363134
rect 37826 327218 38062 327454
rect 38146 327218 38382 327454
rect 37826 326898 38062 327134
rect 38146 326898 38382 327134
rect 37826 291218 38062 291454
rect 38146 291218 38382 291454
rect 37826 290898 38062 291134
rect 38146 290898 38382 291134
rect 37826 255218 38062 255454
rect 38146 255218 38382 255454
rect 37826 254898 38062 255134
rect 38146 254898 38382 255134
rect 37826 219218 38062 219454
rect 38146 219218 38382 219454
rect 37826 218898 38062 219134
rect 38146 218898 38382 219134
rect 37826 183218 38062 183454
rect 38146 183218 38382 183454
rect 37826 182898 38062 183134
rect 38146 182898 38382 183134
rect 37826 147218 38062 147454
rect 38146 147218 38382 147454
rect 37826 146898 38062 147134
rect 38146 146898 38382 147134
rect 37826 111218 38062 111454
rect 38146 111218 38382 111454
rect 37826 110898 38062 111134
rect 38146 110898 38382 111134
rect 37826 75218 38062 75454
rect 38146 75218 38382 75454
rect 37826 74898 38062 75134
rect 38146 74898 38382 75134
rect 37826 39218 38062 39454
rect 38146 39218 38382 39454
rect 37826 38898 38062 39134
rect 38146 38898 38382 39134
rect 37826 3218 38062 3454
rect 38146 3218 38382 3454
rect 37826 2898 38062 3134
rect 38146 2898 38382 3134
rect 37826 -582 38062 -346
rect 38146 -582 38382 -346
rect 37826 -902 38062 -666
rect 38146 -902 38382 -666
rect 41546 690938 41782 691174
rect 41866 690938 42102 691174
rect 41546 690618 41782 690854
rect 41866 690618 42102 690854
rect 41546 654938 41782 655174
rect 41866 654938 42102 655174
rect 41546 654618 41782 654854
rect 41866 654618 42102 654854
rect 41546 618938 41782 619174
rect 41866 618938 42102 619174
rect 41546 618618 41782 618854
rect 41866 618618 42102 618854
rect 41546 582938 41782 583174
rect 41866 582938 42102 583174
rect 41546 582618 41782 582854
rect 41866 582618 42102 582854
rect 41546 546938 41782 547174
rect 41866 546938 42102 547174
rect 41546 546618 41782 546854
rect 41866 546618 42102 546854
rect 41546 510938 41782 511174
rect 41866 510938 42102 511174
rect 41546 510618 41782 510854
rect 41866 510618 42102 510854
rect 41546 474938 41782 475174
rect 41866 474938 42102 475174
rect 41546 474618 41782 474854
rect 41866 474618 42102 474854
rect 41546 438938 41782 439174
rect 41866 438938 42102 439174
rect 41546 438618 41782 438854
rect 41866 438618 42102 438854
rect 41546 402938 41782 403174
rect 41866 402938 42102 403174
rect 41546 402618 41782 402854
rect 41866 402618 42102 402854
rect 41546 366938 41782 367174
rect 41866 366938 42102 367174
rect 41546 366618 41782 366854
rect 41866 366618 42102 366854
rect 41546 330938 41782 331174
rect 41866 330938 42102 331174
rect 41546 330618 41782 330854
rect 41866 330618 42102 330854
rect 41546 294938 41782 295174
rect 41866 294938 42102 295174
rect 41546 294618 41782 294854
rect 41866 294618 42102 294854
rect 41546 258938 41782 259174
rect 41866 258938 42102 259174
rect 41546 258618 41782 258854
rect 41866 258618 42102 258854
rect 41546 222938 41782 223174
rect 41866 222938 42102 223174
rect 41546 222618 41782 222854
rect 41866 222618 42102 222854
rect 41546 186938 41782 187174
rect 41866 186938 42102 187174
rect 41546 186618 41782 186854
rect 41866 186618 42102 186854
rect 41546 150938 41782 151174
rect 41866 150938 42102 151174
rect 41546 150618 41782 150854
rect 41866 150618 42102 150854
rect 41546 114938 41782 115174
rect 41866 114938 42102 115174
rect 41546 114618 41782 114854
rect 41866 114618 42102 114854
rect 41546 78938 41782 79174
rect 41866 78938 42102 79174
rect 41546 78618 41782 78854
rect 41866 78618 42102 78854
rect 41546 42938 41782 43174
rect 41866 42938 42102 43174
rect 41546 42618 41782 42854
rect 41866 42618 42102 42854
rect 41546 6938 41782 7174
rect 41866 6938 42102 7174
rect 41546 6618 41782 6854
rect 41866 6618 42102 6854
rect 41546 -2502 41782 -2266
rect 41866 -2502 42102 -2266
rect 41546 -2822 41782 -2586
rect 41866 -2822 42102 -2586
rect 45266 694658 45502 694894
rect 45586 694658 45822 694894
rect 45266 694338 45502 694574
rect 45586 694338 45822 694574
rect 45266 658658 45502 658894
rect 45586 658658 45822 658894
rect 45266 658338 45502 658574
rect 45586 658338 45822 658574
rect 45266 622658 45502 622894
rect 45586 622658 45822 622894
rect 45266 622338 45502 622574
rect 45586 622338 45822 622574
rect 45266 586658 45502 586894
rect 45586 586658 45822 586894
rect 45266 586338 45502 586574
rect 45586 586338 45822 586574
rect 45266 550658 45502 550894
rect 45586 550658 45822 550894
rect 45266 550338 45502 550574
rect 45586 550338 45822 550574
rect 45266 514658 45502 514894
rect 45586 514658 45822 514894
rect 45266 514338 45502 514574
rect 45586 514338 45822 514574
rect 45266 478658 45502 478894
rect 45586 478658 45822 478894
rect 45266 478338 45502 478574
rect 45586 478338 45822 478574
rect 45266 442658 45502 442894
rect 45586 442658 45822 442894
rect 45266 442338 45502 442574
rect 45586 442338 45822 442574
rect 45266 406658 45502 406894
rect 45586 406658 45822 406894
rect 45266 406338 45502 406574
rect 45586 406338 45822 406574
rect 45266 370658 45502 370894
rect 45586 370658 45822 370894
rect 45266 370338 45502 370574
rect 45586 370338 45822 370574
rect 45266 334658 45502 334894
rect 45586 334658 45822 334894
rect 45266 334338 45502 334574
rect 45586 334338 45822 334574
rect 45266 298658 45502 298894
rect 45586 298658 45822 298894
rect 45266 298338 45502 298574
rect 45586 298338 45822 298574
rect 45266 262658 45502 262894
rect 45586 262658 45822 262894
rect 45266 262338 45502 262574
rect 45586 262338 45822 262574
rect 45266 226658 45502 226894
rect 45586 226658 45822 226894
rect 45266 226338 45502 226574
rect 45586 226338 45822 226574
rect 45266 190658 45502 190894
rect 45586 190658 45822 190894
rect 45266 190338 45502 190574
rect 45586 190338 45822 190574
rect 45266 154658 45502 154894
rect 45586 154658 45822 154894
rect 45266 154338 45502 154574
rect 45586 154338 45822 154574
rect 45266 118658 45502 118894
rect 45586 118658 45822 118894
rect 45266 118338 45502 118574
rect 45586 118338 45822 118574
rect 45266 82658 45502 82894
rect 45586 82658 45822 82894
rect 45266 82338 45502 82574
rect 45586 82338 45822 82574
rect 45266 46658 45502 46894
rect 45586 46658 45822 46894
rect 45266 46338 45502 46574
rect 45586 46338 45822 46574
rect 45266 10658 45502 10894
rect 45586 10658 45822 10894
rect 45266 10338 45502 10574
rect 45586 10338 45822 10574
rect 45266 -4422 45502 -4186
rect 45586 -4422 45822 -4186
rect 45266 -4742 45502 -4506
rect 45586 -4742 45822 -4506
rect 66986 711322 67222 711558
rect 67306 711322 67542 711558
rect 66986 711002 67222 711238
rect 67306 711002 67542 711238
rect 63266 709402 63502 709638
rect 63586 709402 63822 709638
rect 63266 709082 63502 709318
rect 63586 709082 63822 709318
rect 59546 707482 59782 707718
rect 59866 707482 60102 707718
rect 59546 707162 59782 707398
rect 59866 707162 60102 707398
rect 48986 698378 49222 698614
rect 49306 698378 49542 698614
rect 48986 698058 49222 698294
rect 49306 698058 49542 698294
rect 48986 662378 49222 662614
rect 49306 662378 49542 662614
rect 48986 662058 49222 662294
rect 49306 662058 49542 662294
rect 48986 626378 49222 626614
rect 49306 626378 49542 626614
rect 48986 626058 49222 626294
rect 49306 626058 49542 626294
rect 48986 590378 49222 590614
rect 49306 590378 49542 590614
rect 48986 590058 49222 590294
rect 49306 590058 49542 590294
rect 48986 554378 49222 554614
rect 49306 554378 49542 554614
rect 48986 554058 49222 554294
rect 49306 554058 49542 554294
rect 48986 518378 49222 518614
rect 49306 518378 49542 518614
rect 48986 518058 49222 518294
rect 49306 518058 49542 518294
rect 48986 482378 49222 482614
rect 49306 482378 49542 482614
rect 48986 482058 49222 482294
rect 49306 482058 49542 482294
rect 48986 446378 49222 446614
rect 49306 446378 49542 446614
rect 48986 446058 49222 446294
rect 49306 446058 49542 446294
rect 48986 410378 49222 410614
rect 49306 410378 49542 410614
rect 48986 410058 49222 410294
rect 49306 410058 49542 410294
rect 48986 374378 49222 374614
rect 49306 374378 49542 374614
rect 48986 374058 49222 374294
rect 49306 374058 49542 374294
rect 48986 338378 49222 338614
rect 49306 338378 49542 338614
rect 48986 338058 49222 338294
rect 49306 338058 49542 338294
rect 48986 302378 49222 302614
rect 49306 302378 49542 302614
rect 48986 302058 49222 302294
rect 49306 302058 49542 302294
rect 48986 266378 49222 266614
rect 49306 266378 49542 266614
rect 48986 266058 49222 266294
rect 49306 266058 49542 266294
rect 48986 230378 49222 230614
rect 49306 230378 49542 230614
rect 48986 230058 49222 230294
rect 49306 230058 49542 230294
rect 48986 194378 49222 194614
rect 49306 194378 49542 194614
rect 48986 194058 49222 194294
rect 49306 194058 49542 194294
rect 48986 158378 49222 158614
rect 49306 158378 49542 158614
rect 48986 158058 49222 158294
rect 49306 158058 49542 158294
rect 48986 122378 49222 122614
rect 49306 122378 49542 122614
rect 48986 122058 49222 122294
rect 49306 122058 49542 122294
rect 48986 86378 49222 86614
rect 49306 86378 49542 86614
rect 48986 86058 49222 86294
rect 49306 86058 49542 86294
rect 48986 50378 49222 50614
rect 49306 50378 49542 50614
rect 48986 50058 49222 50294
rect 49306 50058 49542 50294
rect 48986 14378 49222 14614
rect 49306 14378 49542 14614
rect 48986 14058 49222 14294
rect 49306 14058 49542 14294
rect 30986 -7302 31222 -7066
rect 31306 -7302 31542 -7066
rect 30986 -7622 31222 -7386
rect 31306 -7622 31542 -7386
rect 55826 705562 56062 705798
rect 56146 705562 56382 705798
rect 55826 705242 56062 705478
rect 56146 705242 56382 705478
rect 55826 669218 56062 669454
rect 56146 669218 56382 669454
rect 55826 668898 56062 669134
rect 56146 668898 56382 669134
rect 55826 633218 56062 633454
rect 56146 633218 56382 633454
rect 55826 632898 56062 633134
rect 56146 632898 56382 633134
rect 55826 597218 56062 597454
rect 56146 597218 56382 597454
rect 55826 596898 56062 597134
rect 56146 596898 56382 597134
rect 55826 561218 56062 561454
rect 56146 561218 56382 561454
rect 55826 560898 56062 561134
rect 56146 560898 56382 561134
rect 55826 525218 56062 525454
rect 56146 525218 56382 525454
rect 55826 524898 56062 525134
rect 56146 524898 56382 525134
rect 55826 489218 56062 489454
rect 56146 489218 56382 489454
rect 55826 488898 56062 489134
rect 56146 488898 56382 489134
rect 55826 453218 56062 453454
rect 56146 453218 56382 453454
rect 55826 452898 56062 453134
rect 56146 452898 56382 453134
rect 55826 417218 56062 417454
rect 56146 417218 56382 417454
rect 55826 416898 56062 417134
rect 56146 416898 56382 417134
rect 55826 381218 56062 381454
rect 56146 381218 56382 381454
rect 55826 380898 56062 381134
rect 56146 380898 56382 381134
rect 55826 345218 56062 345454
rect 56146 345218 56382 345454
rect 55826 344898 56062 345134
rect 56146 344898 56382 345134
rect 55826 309218 56062 309454
rect 56146 309218 56382 309454
rect 55826 308898 56062 309134
rect 56146 308898 56382 309134
rect 55826 273218 56062 273454
rect 56146 273218 56382 273454
rect 55826 272898 56062 273134
rect 56146 272898 56382 273134
rect 55826 237218 56062 237454
rect 56146 237218 56382 237454
rect 55826 236898 56062 237134
rect 56146 236898 56382 237134
rect 55826 201218 56062 201454
rect 56146 201218 56382 201454
rect 55826 200898 56062 201134
rect 56146 200898 56382 201134
rect 55826 165218 56062 165454
rect 56146 165218 56382 165454
rect 55826 164898 56062 165134
rect 56146 164898 56382 165134
rect 55826 129218 56062 129454
rect 56146 129218 56382 129454
rect 55826 128898 56062 129134
rect 56146 128898 56382 129134
rect 55826 93218 56062 93454
rect 56146 93218 56382 93454
rect 55826 92898 56062 93134
rect 56146 92898 56382 93134
rect 55826 57218 56062 57454
rect 56146 57218 56382 57454
rect 55826 56898 56062 57134
rect 56146 56898 56382 57134
rect 55826 21218 56062 21454
rect 56146 21218 56382 21454
rect 55826 20898 56062 21134
rect 56146 20898 56382 21134
rect 55826 -1542 56062 -1306
rect 56146 -1542 56382 -1306
rect 55826 -1862 56062 -1626
rect 56146 -1862 56382 -1626
rect 59546 672938 59782 673174
rect 59866 672938 60102 673174
rect 59546 672618 59782 672854
rect 59866 672618 60102 672854
rect 59546 636938 59782 637174
rect 59866 636938 60102 637174
rect 59546 636618 59782 636854
rect 59866 636618 60102 636854
rect 59546 600938 59782 601174
rect 59866 600938 60102 601174
rect 59546 600618 59782 600854
rect 59866 600618 60102 600854
rect 59546 564938 59782 565174
rect 59866 564938 60102 565174
rect 59546 564618 59782 564854
rect 59866 564618 60102 564854
rect 59546 528938 59782 529174
rect 59866 528938 60102 529174
rect 59546 528618 59782 528854
rect 59866 528618 60102 528854
rect 59546 492938 59782 493174
rect 59866 492938 60102 493174
rect 59546 492618 59782 492854
rect 59866 492618 60102 492854
rect 59546 456938 59782 457174
rect 59866 456938 60102 457174
rect 59546 456618 59782 456854
rect 59866 456618 60102 456854
rect 59546 420938 59782 421174
rect 59866 420938 60102 421174
rect 59546 420618 59782 420854
rect 59866 420618 60102 420854
rect 59546 384938 59782 385174
rect 59866 384938 60102 385174
rect 59546 384618 59782 384854
rect 59866 384618 60102 384854
rect 59546 348938 59782 349174
rect 59866 348938 60102 349174
rect 59546 348618 59782 348854
rect 59866 348618 60102 348854
rect 59546 312938 59782 313174
rect 59866 312938 60102 313174
rect 59546 312618 59782 312854
rect 59866 312618 60102 312854
rect 59546 276938 59782 277174
rect 59866 276938 60102 277174
rect 59546 276618 59782 276854
rect 59866 276618 60102 276854
rect 59546 240938 59782 241174
rect 59866 240938 60102 241174
rect 59546 240618 59782 240854
rect 59866 240618 60102 240854
rect 59546 204938 59782 205174
rect 59866 204938 60102 205174
rect 59546 204618 59782 204854
rect 59866 204618 60102 204854
rect 59546 168938 59782 169174
rect 59866 168938 60102 169174
rect 59546 168618 59782 168854
rect 59866 168618 60102 168854
rect 59546 132938 59782 133174
rect 59866 132938 60102 133174
rect 59546 132618 59782 132854
rect 59866 132618 60102 132854
rect 59546 96938 59782 97174
rect 59866 96938 60102 97174
rect 59546 96618 59782 96854
rect 59866 96618 60102 96854
rect 59546 60938 59782 61174
rect 59866 60938 60102 61174
rect 59546 60618 59782 60854
rect 59866 60618 60102 60854
rect 59546 24938 59782 25174
rect 59866 24938 60102 25174
rect 59546 24618 59782 24854
rect 59866 24618 60102 24854
rect 59546 -3462 59782 -3226
rect 59866 -3462 60102 -3226
rect 59546 -3782 59782 -3546
rect 59866 -3782 60102 -3546
rect 63266 676658 63502 676894
rect 63586 676658 63822 676894
rect 63266 676338 63502 676574
rect 63586 676338 63822 676574
rect 63266 640658 63502 640894
rect 63586 640658 63822 640894
rect 63266 640338 63502 640574
rect 63586 640338 63822 640574
rect 63266 604658 63502 604894
rect 63586 604658 63822 604894
rect 63266 604338 63502 604574
rect 63586 604338 63822 604574
rect 63266 568658 63502 568894
rect 63586 568658 63822 568894
rect 63266 568338 63502 568574
rect 63586 568338 63822 568574
rect 63266 532658 63502 532894
rect 63586 532658 63822 532894
rect 63266 532338 63502 532574
rect 63586 532338 63822 532574
rect 63266 496658 63502 496894
rect 63586 496658 63822 496894
rect 63266 496338 63502 496574
rect 63586 496338 63822 496574
rect 63266 460658 63502 460894
rect 63586 460658 63822 460894
rect 63266 460338 63502 460574
rect 63586 460338 63822 460574
rect 63266 424658 63502 424894
rect 63586 424658 63822 424894
rect 63266 424338 63502 424574
rect 63586 424338 63822 424574
rect 63266 388658 63502 388894
rect 63586 388658 63822 388894
rect 63266 388338 63502 388574
rect 63586 388338 63822 388574
rect 63266 352658 63502 352894
rect 63586 352658 63822 352894
rect 63266 352338 63502 352574
rect 63586 352338 63822 352574
rect 63266 316658 63502 316894
rect 63586 316658 63822 316894
rect 63266 316338 63502 316574
rect 63586 316338 63822 316574
rect 63266 280658 63502 280894
rect 63586 280658 63822 280894
rect 63266 280338 63502 280574
rect 63586 280338 63822 280574
rect 63266 244658 63502 244894
rect 63586 244658 63822 244894
rect 63266 244338 63502 244574
rect 63586 244338 63822 244574
rect 63266 208658 63502 208894
rect 63586 208658 63822 208894
rect 63266 208338 63502 208574
rect 63586 208338 63822 208574
rect 63266 172658 63502 172894
rect 63586 172658 63822 172894
rect 63266 172338 63502 172574
rect 63586 172338 63822 172574
rect 63266 136658 63502 136894
rect 63586 136658 63822 136894
rect 63266 136338 63502 136574
rect 63586 136338 63822 136574
rect 63266 100658 63502 100894
rect 63586 100658 63822 100894
rect 63266 100338 63502 100574
rect 63586 100338 63822 100574
rect 63266 64658 63502 64894
rect 63586 64658 63822 64894
rect 63266 64338 63502 64574
rect 63586 64338 63822 64574
rect 63266 28658 63502 28894
rect 63586 28658 63822 28894
rect 63266 28338 63502 28574
rect 63586 28338 63822 28574
rect 63266 -5382 63502 -5146
rect 63586 -5382 63822 -5146
rect 63266 -5702 63502 -5466
rect 63586 -5702 63822 -5466
rect 84986 710362 85222 710598
rect 85306 710362 85542 710598
rect 84986 710042 85222 710278
rect 85306 710042 85542 710278
rect 81266 708442 81502 708678
rect 81586 708442 81822 708678
rect 81266 708122 81502 708358
rect 81586 708122 81822 708358
rect 77546 706522 77782 706758
rect 77866 706522 78102 706758
rect 77546 706202 77782 706438
rect 77866 706202 78102 706438
rect 66986 680378 67222 680614
rect 67306 680378 67542 680614
rect 66986 680058 67222 680294
rect 67306 680058 67542 680294
rect 66986 644378 67222 644614
rect 67306 644378 67542 644614
rect 66986 644058 67222 644294
rect 67306 644058 67542 644294
rect 66986 608378 67222 608614
rect 67306 608378 67542 608614
rect 66986 608058 67222 608294
rect 67306 608058 67542 608294
rect 66986 572378 67222 572614
rect 67306 572378 67542 572614
rect 66986 572058 67222 572294
rect 67306 572058 67542 572294
rect 66986 536378 67222 536614
rect 67306 536378 67542 536614
rect 66986 536058 67222 536294
rect 67306 536058 67542 536294
rect 66986 500378 67222 500614
rect 67306 500378 67542 500614
rect 66986 500058 67222 500294
rect 67306 500058 67542 500294
rect 66986 464378 67222 464614
rect 67306 464378 67542 464614
rect 66986 464058 67222 464294
rect 67306 464058 67542 464294
rect 66986 428378 67222 428614
rect 67306 428378 67542 428614
rect 66986 428058 67222 428294
rect 67306 428058 67542 428294
rect 66986 392378 67222 392614
rect 67306 392378 67542 392614
rect 66986 392058 67222 392294
rect 67306 392058 67542 392294
rect 66986 356378 67222 356614
rect 67306 356378 67542 356614
rect 66986 356058 67222 356294
rect 67306 356058 67542 356294
rect 66986 320378 67222 320614
rect 67306 320378 67542 320614
rect 66986 320058 67222 320294
rect 67306 320058 67542 320294
rect 66986 284378 67222 284614
rect 67306 284378 67542 284614
rect 66986 284058 67222 284294
rect 67306 284058 67542 284294
rect 66986 248378 67222 248614
rect 67306 248378 67542 248614
rect 66986 248058 67222 248294
rect 67306 248058 67542 248294
rect 66986 212378 67222 212614
rect 67306 212378 67542 212614
rect 66986 212058 67222 212294
rect 67306 212058 67542 212294
rect 66986 176378 67222 176614
rect 67306 176378 67542 176614
rect 66986 176058 67222 176294
rect 67306 176058 67542 176294
rect 66986 140378 67222 140614
rect 67306 140378 67542 140614
rect 66986 140058 67222 140294
rect 67306 140058 67542 140294
rect 66986 104378 67222 104614
rect 67306 104378 67542 104614
rect 66986 104058 67222 104294
rect 67306 104058 67542 104294
rect 66986 68378 67222 68614
rect 67306 68378 67542 68614
rect 66986 68058 67222 68294
rect 67306 68058 67542 68294
rect 66986 32378 67222 32614
rect 67306 32378 67542 32614
rect 66986 32058 67222 32294
rect 67306 32058 67542 32294
rect 48986 -6342 49222 -6106
rect 49306 -6342 49542 -6106
rect 48986 -6662 49222 -6426
rect 49306 -6662 49542 -6426
rect 73826 704602 74062 704838
rect 74146 704602 74382 704838
rect 73826 704282 74062 704518
rect 74146 704282 74382 704518
rect 73826 687218 74062 687454
rect 74146 687218 74382 687454
rect 73826 686898 74062 687134
rect 74146 686898 74382 687134
rect 73826 651218 74062 651454
rect 74146 651218 74382 651454
rect 73826 650898 74062 651134
rect 74146 650898 74382 651134
rect 73826 615218 74062 615454
rect 74146 615218 74382 615454
rect 73826 614898 74062 615134
rect 74146 614898 74382 615134
rect 73826 579218 74062 579454
rect 74146 579218 74382 579454
rect 73826 578898 74062 579134
rect 74146 578898 74382 579134
rect 73826 543218 74062 543454
rect 74146 543218 74382 543454
rect 73826 542898 74062 543134
rect 74146 542898 74382 543134
rect 73826 507218 74062 507454
rect 74146 507218 74382 507454
rect 73826 506898 74062 507134
rect 74146 506898 74382 507134
rect 73826 471218 74062 471454
rect 74146 471218 74382 471454
rect 73826 470898 74062 471134
rect 74146 470898 74382 471134
rect 73826 435218 74062 435454
rect 74146 435218 74382 435454
rect 73826 434898 74062 435134
rect 74146 434898 74382 435134
rect 73826 399218 74062 399454
rect 74146 399218 74382 399454
rect 73826 398898 74062 399134
rect 74146 398898 74382 399134
rect 73826 363218 74062 363454
rect 74146 363218 74382 363454
rect 73826 362898 74062 363134
rect 74146 362898 74382 363134
rect 73826 327218 74062 327454
rect 74146 327218 74382 327454
rect 73826 326898 74062 327134
rect 74146 326898 74382 327134
rect 73826 291218 74062 291454
rect 74146 291218 74382 291454
rect 73826 290898 74062 291134
rect 74146 290898 74382 291134
rect 73826 255218 74062 255454
rect 74146 255218 74382 255454
rect 73826 254898 74062 255134
rect 74146 254898 74382 255134
rect 73826 219218 74062 219454
rect 74146 219218 74382 219454
rect 73826 218898 74062 219134
rect 74146 218898 74382 219134
rect 73826 183218 74062 183454
rect 74146 183218 74382 183454
rect 73826 182898 74062 183134
rect 74146 182898 74382 183134
rect 73826 147218 74062 147454
rect 74146 147218 74382 147454
rect 73826 146898 74062 147134
rect 74146 146898 74382 147134
rect 73826 111218 74062 111454
rect 74146 111218 74382 111454
rect 73826 110898 74062 111134
rect 74146 110898 74382 111134
rect 73826 75218 74062 75454
rect 74146 75218 74382 75454
rect 73826 74898 74062 75134
rect 74146 74898 74382 75134
rect 73826 39218 74062 39454
rect 74146 39218 74382 39454
rect 73826 38898 74062 39134
rect 74146 38898 74382 39134
rect 73826 3218 74062 3454
rect 74146 3218 74382 3454
rect 73826 2898 74062 3134
rect 74146 2898 74382 3134
rect 73826 -582 74062 -346
rect 74146 -582 74382 -346
rect 73826 -902 74062 -666
rect 74146 -902 74382 -666
rect 77546 690938 77782 691174
rect 77866 690938 78102 691174
rect 77546 690618 77782 690854
rect 77866 690618 78102 690854
rect 77546 654938 77782 655174
rect 77866 654938 78102 655174
rect 77546 654618 77782 654854
rect 77866 654618 78102 654854
rect 77546 618938 77782 619174
rect 77866 618938 78102 619174
rect 77546 618618 77782 618854
rect 77866 618618 78102 618854
rect 77546 582938 77782 583174
rect 77866 582938 78102 583174
rect 77546 582618 77782 582854
rect 77866 582618 78102 582854
rect 77546 546938 77782 547174
rect 77866 546938 78102 547174
rect 77546 546618 77782 546854
rect 77866 546618 78102 546854
rect 77546 510938 77782 511174
rect 77866 510938 78102 511174
rect 77546 510618 77782 510854
rect 77866 510618 78102 510854
rect 77546 474938 77782 475174
rect 77866 474938 78102 475174
rect 77546 474618 77782 474854
rect 77866 474618 78102 474854
rect 77546 438938 77782 439174
rect 77866 438938 78102 439174
rect 77546 438618 77782 438854
rect 77866 438618 78102 438854
rect 77546 402938 77782 403174
rect 77866 402938 78102 403174
rect 77546 402618 77782 402854
rect 77866 402618 78102 402854
rect 77546 366938 77782 367174
rect 77866 366938 78102 367174
rect 77546 366618 77782 366854
rect 77866 366618 78102 366854
rect 77546 330938 77782 331174
rect 77866 330938 78102 331174
rect 77546 330618 77782 330854
rect 77866 330618 78102 330854
rect 77546 294938 77782 295174
rect 77866 294938 78102 295174
rect 77546 294618 77782 294854
rect 77866 294618 78102 294854
rect 77546 258938 77782 259174
rect 77866 258938 78102 259174
rect 77546 258618 77782 258854
rect 77866 258618 78102 258854
rect 77546 222938 77782 223174
rect 77866 222938 78102 223174
rect 77546 222618 77782 222854
rect 77866 222618 78102 222854
rect 77546 186938 77782 187174
rect 77866 186938 78102 187174
rect 77546 186618 77782 186854
rect 77866 186618 78102 186854
rect 77546 150938 77782 151174
rect 77866 150938 78102 151174
rect 77546 150618 77782 150854
rect 77866 150618 78102 150854
rect 77546 114938 77782 115174
rect 77866 114938 78102 115174
rect 77546 114618 77782 114854
rect 77866 114618 78102 114854
rect 77546 78938 77782 79174
rect 77866 78938 78102 79174
rect 77546 78618 77782 78854
rect 77866 78618 78102 78854
rect 77546 42938 77782 43174
rect 77866 42938 78102 43174
rect 77546 42618 77782 42854
rect 77866 42618 78102 42854
rect 77546 6938 77782 7174
rect 77866 6938 78102 7174
rect 77546 6618 77782 6854
rect 77866 6618 78102 6854
rect 77546 -2502 77782 -2266
rect 77866 -2502 78102 -2266
rect 77546 -2822 77782 -2586
rect 77866 -2822 78102 -2586
rect 81266 694658 81502 694894
rect 81586 694658 81822 694894
rect 81266 694338 81502 694574
rect 81586 694338 81822 694574
rect 81266 658658 81502 658894
rect 81586 658658 81822 658894
rect 81266 658338 81502 658574
rect 81586 658338 81822 658574
rect 81266 622658 81502 622894
rect 81586 622658 81822 622894
rect 81266 622338 81502 622574
rect 81586 622338 81822 622574
rect 81266 586658 81502 586894
rect 81586 586658 81822 586894
rect 81266 586338 81502 586574
rect 81586 586338 81822 586574
rect 81266 550658 81502 550894
rect 81586 550658 81822 550894
rect 81266 550338 81502 550574
rect 81586 550338 81822 550574
rect 81266 514658 81502 514894
rect 81586 514658 81822 514894
rect 81266 514338 81502 514574
rect 81586 514338 81822 514574
rect 81266 478658 81502 478894
rect 81586 478658 81822 478894
rect 81266 478338 81502 478574
rect 81586 478338 81822 478574
rect 81266 442658 81502 442894
rect 81586 442658 81822 442894
rect 81266 442338 81502 442574
rect 81586 442338 81822 442574
rect 81266 406658 81502 406894
rect 81586 406658 81822 406894
rect 81266 406338 81502 406574
rect 81586 406338 81822 406574
rect 81266 370658 81502 370894
rect 81586 370658 81822 370894
rect 81266 370338 81502 370574
rect 81586 370338 81822 370574
rect 81266 334658 81502 334894
rect 81586 334658 81822 334894
rect 81266 334338 81502 334574
rect 81586 334338 81822 334574
rect 81266 298658 81502 298894
rect 81586 298658 81822 298894
rect 81266 298338 81502 298574
rect 81586 298338 81822 298574
rect 81266 262658 81502 262894
rect 81586 262658 81822 262894
rect 81266 262338 81502 262574
rect 81586 262338 81822 262574
rect 81266 226658 81502 226894
rect 81586 226658 81822 226894
rect 81266 226338 81502 226574
rect 81586 226338 81822 226574
rect 81266 190658 81502 190894
rect 81586 190658 81822 190894
rect 81266 190338 81502 190574
rect 81586 190338 81822 190574
rect 81266 154658 81502 154894
rect 81586 154658 81822 154894
rect 81266 154338 81502 154574
rect 81586 154338 81822 154574
rect 81266 118658 81502 118894
rect 81586 118658 81822 118894
rect 81266 118338 81502 118574
rect 81586 118338 81822 118574
rect 81266 82658 81502 82894
rect 81586 82658 81822 82894
rect 81266 82338 81502 82574
rect 81586 82338 81822 82574
rect 81266 46658 81502 46894
rect 81586 46658 81822 46894
rect 81266 46338 81502 46574
rect 81586 46338 81822 46574
rect 81266 10658 81502 10894
rect 81586 10658 81822 10894
rect 81266 10338 81502 10574
rect 81586 10338 81822 10574
rect 81266 -4422 81502 -4186
rect 81586 -4422 81822 -4186
rect 81266 -4742 81502 -4506
rect 81586 -4742 81822 -4506
rect 102986 711322 103222 711558
rect 103306 711322 103542 711558
rect 102986 711002 103222 711238
rect 103306 711002 103542 711238
rect 99266 709402 99502 709638
rect 99586 709402 99822 709638
rect 99266 709082 99502 709318
rect 99586 709082 99822 709318
rect 95546 707482 95782 707718
rect 95866 707482 96102 707718
rect 95546 707162 95782 707398
rect 95866 707162 96102 707398
rect 84986 698378 85222 698614
rect 85306 698378 85542 698614
rect 84986 698058 85222 698294
rect 85306 698058 85542 698294
rect 84986 662378 85222 662614
rect 85306 662378 85542 662614
rect 84986 662058 85222 662294
rect 85306 662058 85542 662294
rect 84986 626378 85222 626614
rect 85306 626378 85542 626614
rect 84986 626058 85222 626294
rect 85306 626058 85542 626294
rect 84986 590378 85222 590614
rect 85306 590378 85542 590614
rect 84986 590058 85222 590294
rect 85306 590058 85542 590294
rect 84986 554378 85222 554614
rect 85306 554378 85542 554614
rect 84986 554058 85222 554294
rect 85306 554058 85542 554294
rect 84986 518378 85222 518614
rect 85306 518378 85542 518614
rect 84986 518058 85222 518294
rect 85306 518058 85542 518294
rect 84986 482378 85222 482614
rect 85306 482378 85542 482614
rect 84986 482058 85222 482294
rect 85306 482058 85542 482294
rect 84986 446378 85222 446614
rect 85306 446378 85542 446614
rect 84986 446058 85222 446294
rect 85306 446058 85542 446294
rect 84986 410378 85222 410614
rect 85306 410378 85542 410614
rect 84986 410058 85222 410294
rect 85306 410058 85542 410294
rect 84986 374378 85222 374614
rect 85306 374378 85542 374614
rect 84986 374058 85222 374294
rect 85306 374058 85542 374294
rect 84986 338378 85222 338614
rect 85306 338378 85542 338614
rect 84986 338058 85222 338294
rect 85306 338058 85542 338294
rect 84986 302378 85222 302614
rect 85306 302378 85542 302614
rect 84986 302058 85222 302294
rect 85306 302058 85542 302294
rect 84986 266378 85222 266614
rect 85306 266378 85542 266614
rect 84986 266058 85222 266294
rect 85306 266058 85542 266294
rect 84986 230378 85222 230614
rect 85306 230378 85542 230614
rect 84986 230058 85222 230294
rect 85306 230058 85542 230294
rect 84986 194378 85222 194614
rect 85306 194378 85542 194614
rect 84986 194058 85222 194294
rect 85306 194058 85542 194294
rect 84986 158378 85222 158614
rect 85306 158378 85542 158614
rect 84986 158058 85222 158294
rect 85306 158058 85542 158294
rect 84986 122378 85222 122614
rect 85306 122378 85542 122614
rect 84986 122058 85222 122294
rect 85306 122058 85542 122294
rect 84986 86378 85222 86614
rect 85306 86378 85542 86614
rect 84986 86058 85222 86294
rect 85306 86058 85542 86294
rect 84986 50378 85222 50614
rect 85306 50378 85542 50614
rect 84986 50058 85222 50294
rect 85306 50058 85542 50294
rect 84986 14378 85222 14614
rect 85306 14378 85542 14614
rect 84986 14058 85222 14294
rect 85306 14058 85542 14294
rect 66986 -7302 67222 -7066
rect 67306 -7302 67542 -7066
rect 66986 -7622 67222 -7386
rect 67306 -7622 67542 -7386
rect 91826 705562 92062 705798
rect 92146 705562 92382 705798
rect 91826 705242 92062 705478
rect 92146 705242 92382 705478
rect 91826 669218 92062 669454
rect 92146 669218 92382 669454
rect 91826 668898 92062 669134
rect 92146 668898 92382 669134
rect 91826 633218 92062 633454
rect 92146 633218 92382 633454
rect 91826 632898 92062 633134
rect 92146 632898 92382 633134
rect 91826 597218 92062 597454
rect 92146 597218 92382 597454
rect 91826 596898 92062 597134
rect 92146 596898 92382 597134
rect 91826 561218 92062 561454
rect 92146 561218 92382 561454
rect 91826 560898 92062 561134
rect 92146 560898 92382 561134
rect 91826 525218 92062 525454
rect 92146 525218 92382 525454
rect 91826 524898 92062 525134
rect 92146 524898 92382 525134
rect 91826 489218 92062 489454
rect 92146 489218 92382 489454
rect 91826 488898 92062 489134
rect 92146 488898 92382 489134
rect 91826 453218 92062 453454
rect 92146 453218 92382 453454
rect 91826 452898 92062 453134
rect 92146 452898 92382 453134
rect 91826 417218 92062 417454
rect 92146 417218 92382 417454
rect 91826 416898 92062 417134
rect 92146 416898 92382 417134
rect 91826 381218 92062 381454
rect 92146 381218 92382 381454
rect 91826 380898 92062 381134
rect 92146 380898 92382 381134
rect 91826 345218 92062 345454
rect 92146 345218 92382 345454
rect 91826 344898 92062 345134
rect 92146 344898 92382 345134
rect 91826 309218 92062 309454
rect 92146 309218 92382 309454
rect 91826 308898 92062 309134
rect 92146 308898 92382 309134
rect 91826 273218 92062 273454
rect 92146 273218 92382 273454
rect 91826 272898 92062 273134
rect 92146 272898 92382 273134
rect 91826 237218 92062 237454
rect 92146 237218 92382 237454
rect 91826 236898 92062 237134
rect 92146 236898 92382 237134
rect 91826 201218 92062 201454
rect 92146 201218 92382 201454
rect 91826 200898 92062 201134
rect 92146 200898 92382 201134
rect 91826 165218 92062 165454
rect 92146 165218 92382 165454
rect 91826 164898 92062 165134
rect 92146 164898 92382 165134
rect 91826 129218 92062 129454
rect 92146 129218 92382 129454
rect 91826 128898 92062 129134
rect 92146 128898 92382 129134
rect 91826 93218 92062 93454
rect 92146 93218 92382 93454
rect 91826 92898 92062 93134
rect 92146 92898 92382 93134
rect 91826 57218 92062 57454
rect 92146 57218 92382 57454
rect 91826 56898 92062 57134
rect 92146 56898 92382 57134
rect 91826 21218 92062 21454
rect 92146 21218 92382 21454
rect 91826 20898 92062 21134
rect 92146 20898 92382 21134
rect 91826 -1542 92062 -1306
rect 92146 -1542 92382 -1306
rect 91826 -1862 92062 -1626
rect 92146 -1862 92382 -1626
rect 95546 672938 95782 673174
rect 95866 672938 96102 673174
rect 95546 672618 95782 672854
rect 95866 672618 96102 672854
rect 95546 636938 95782 637174
rect 95866 636938 96102 637174
rect 95546 636618 95782 636854
rect 95866 636618 96102 636854
rect 95546 600938 95782 601174
rect 95866 600938 96102 601174
rect 95546 600618 95782 600854
rect 95866 600618 96102 600854
rect 95546 564938 95782 565174
rect 95866 564938 96102 565174
rect 95546 564618 95782 564854
rect 95866 564618 96102 564854
rect 95546 528938 95782 529174
rect 95866 528938 96102 529174
rect 95546 528618 95782 528854
rect 95866 528618 96102 528854
rect 95546 492938 95782 493174
rect 95866 492938 96102 493174
rect 95546 492618 95782 492854
rect 95866 492618 96102 492854
rect 95546 456938 95782 457174
rect 95866 456938 96102 457174
rect 95546 456618 95782 456854
rect 95866 456618 96102 456854
rect 95546 420938 95782 421174
rect 95866 420938 96102 421174
rect 95546 420618 95782 420854
rect 95866 420618 96102 420854
rect 95546 384938 95782 385174
rect 95866 384938 96102 385174
rect 95546 384618 95782 384854
rect 95866 384618 96102 384854
rect 95546 348938 95782 349174
rect 95866 348938 96102 349174
rect 95546 348618 95782 348854
rect 95866 348618 96102 348854
rect 95546 312938 95782 313174
rect 95866 312938 96102 313174
rect 95546 312618 95782 312854
rect 95866 312618 96102 312854
rect 95546 276938 95782 277174
rect 95866 276938 96102 277174
rect 95546 276618 95782 276854
rect 95866 276618 96102 276854
rect 95546 240938 95782 241174
rect 95866 240938 96102 241174
rect 95546 240618 95782 240854
rect 95866 240618 96102 240854
rect 95546 204938 95782 205174
rect 95866 204938 96102 205174
rect 95546 204618 95782 204854
rect 95866 204618 96102 204854
rect 95546 168938 95782 169174
rect 95866 168938 96102 169174
rect 95546 168618 95782 168854
rect 95866 168618 96102 168854
rect 95546 132938 95782 133174
rect 95866 132938 96102 133174
rect 95546 132618 95782 132854
rect 95866 132618 96102 132854
rect 95546 96938 95782 97174
rect 95866 96938 96102 97174
rect 95546 96618 95782 96854
rect 95866 96618 96102 96854
rect 95546 60938 95782 61174
rect 95866 60938 96102 61174
rect 95546 60618 95782 60854
rect 95866 60618 96102 60854
rect 95546 24938 95782 25174
rect 95866 24938 96102 25174
rect 95546 24618 95782 24854
rect 95866 24618 96102 24854
rect 95546 -3462 95782 -3226
rect 95866 -3462 96102 -3226
rect 95546 -3782 95782 -3546
rect 95866 -3782 96102 -3546
rect 99266 676658 99502 676894
rect 99586 676658 99822 676894
rect 99266 676338 99502 676574
rect 99586 676338 99822 676574
rect 99266 640658 99502 640894
rect 99586 640658 99822 640894
rect 99266 640338 99502 640574
rect 99586 640338 99822 640574
rect 99266 604658 99502 604894
rect 99586 604658 99822 604894
rect 99266 604338 99502 604574
rect 99586 604338 99822 604574
rect 99266 568658 99502 568894
rect 99586 568658 99822 568894
rect 99266 568338 99502 568574
rect 99586 568338 99822 568574
rect 99266 532658 99502 532894
rect 99586 532658 99822 532894
rect 99266 532338 99502 532574
rect 99586 532338 99822 532574
rect 99266 496658 99502 496894
rect 99586 496658 99822 496894
rect 99266 496338 99502 496574
rect 99586 496338 99822 496574
rect 99266 460658 99502 460894
rect 99586 460658 99822 460894
rect 99266 460338 99502 460574
rect 99586 460338 99822 460574
rect 99266 424658 99502 424894
rect 99586 424658 99822 424894
rect 99266 424338 99502 424574
rect 99586 424338 99822 424574
rect 99266 388658 99502 388894
rect 99586 388658 99822 388894
rect 99266 388338 99502 388574
rect 99586 388338 99822 388574
rect 99266 352658 99502 352894
rect 99586 352658 99822 352894
rect 99266 352338 99502 352574
rect 99586 352338 99822 352574
rect 99266 316658 99502 316894
rect 99586 316658 99822 316894
rect 99266 316338 99502 316574
rect 99586 316338 99822 316574
rect 99266 280658 99502 280894
rect 99586 280658 99822 280894
rect 99266 280338 99502 280574
rect 99586 280338 99822 280574
rect 99266 244658 99502 244894
rect 99586 244658 99822 244894
rect 99266 244338 99502 244574
rect 99586 244338 99822 244574
rect 99266 208658 99502 208894
rect 99586 208658 99822 208894
rect 99266 208338 99502 208574
rect 99586 208338 99822 208574
rect 99266 172658 99502 172894
rect 99586 172658 99822 172894
rect 99266 172338 99502 172574
rect 99586 172338 99822 172574
rect 99266 136658 99502 136894
rect 99586 136658 99822 136894
rect 99266 136338 99502 136574
rect 99586 136338 99822 136574
rect 99266 100658 99502 100894
rect 99586 100658 99822 100894
rect 99266 100338 99502 100574
rect 99586 100338 99822 100574
rect 99266 64658 99502 64894
rect 99586 64658 99822 64894
rect 99266 64338 99502 64574
rect 99586 64338 99822 64574
rect 99266 28658 99502 28894
rect 99586 28658 99822 28894
rect 99266 28338 99502 28574
rect 99586 28338 99822 28574
rect 99266 -5382 99502 -5146
rect 99586 -5382 99822 -5146
rect 99266 -5702 99502 -5466
rect 99586 -5702 99822 -5466
rect 120986 710362 121222 710598
rect 121306 710362 121542 710598
rect 120986 710042 121222 710278
rect 121306 710042 121542 710278
rect 117266 708442 117502 708678
rect 117586 708442 117822 708678
rect 117266 708122 117502 708358
rect 117586 708122 117822 708358
rect 113546 706522 113782 706758
rect 113866 706522 114102 706758
rect 113546 706202 113782 706438
rect 113866 706202 114102 706438
rect 102986 680378 103222 680614
rect 103306 680378 103542 680614
rect 102986 680058 103222 680294
rect 103306 680058 103542 680294
rect 102986 644378 103222 644614
rect 103306 644378 103542 644614
rect 102986 644058 103222 644294
rect 103306 644058 103542 644294
rect 102986 608378 103222 608614
rect 103306 608378 103542 608614
rect 102986 608058 103222 608294
rect 103306 608058 103542 608294
rect 102986 572378 103222 572614
rect 103306 572378 103542 572614
rect 102986 572058 103222 572294
rect 103306 572058 103542 572294
rect 102986 536378 103222 536614
rect 103306 536378 103542 536614
rect 102986 536058 103222 536294
rect 103306 536058 103542 536294
rect 102986 500378 103222 500614
rect 103306 500378 103542 500614
rect 102986 500058 103222 500294
rect 103306 500058 103542 500294
rect 102986 464378 103222 464614
rect 103306 464378 103542 464614
rect 102986 464058 103222 464294
rect 103306 464058 103542 464294
rect 102986 428378 103222 428614
rect 103306 428378 103542 428614
rect 102986 428058 103222 428294
rect 103306 428058 103542 428294
rect 102986 392378 103222 392614
rect 103306 392378 103542 392614
rect 102986 392058 103222 392294
rect 103306 392058 103542 392294
rect 102986 356378 103222 356614
rect 103306 356378 103542 356614
rect 102986 356058 103222 356294
rect 103306 356058 103542 356294
rect 102986 320378 103222 320614
rect 103306 320378 103542 320614
rect 102986 320058 103222 320294
rect 103306 320058 103542 320294
rect 102986 284378 103222 284614
rect 103306 284378 103542 284614
rect 102986 284058 103222 284294
rect 103306 284058 103542 284294
rect 102986 248378 103222 248614
rect 103306 248378 103542 248614
rect 102986 248058 103222 248294
rect 103306 248058 103542 248294
rect 102986 212378 103222 212614
rect 103306 212378 103542 212614
rect 102986 212058 103222 212294
rect 103306 212058 103542 212294
rect 102986 176378 103222 176614
rect 103306 176378 103542 176614
rect 102986 176058 103222 176294
rect 103306 176058 103542 176294
rect 102986 140378 103222 140614
rect 103306 140378 103542 140614
rect 102986 140058 103222 140294
rect 103306 140058 103542 140294
rect 102986 104378 103222 104614
rect 103306 104378 103542 104614
rect 102986 104058 103222 104294
rect 103306 104058 103542 104294
rect 102986 68378 103222 68614
rect 103306 68378 103542 68614
rect 102986 68058 103222 68294
rect 103306 68058 103542 68294
rect 102986 32378 103222 32614
rect 103306 32378 103542 32614
rect 102986 32058 103222 32294
rect 103306 32058 103542 32294
rect 84986 -6342 85222 -6106
rect 85306 -6342 85542 -6106
rect 84986 -6662 85222 -6426
rect 85306 -6662 85542 -6426
rect 109826 704602 110062 704838
rect 110146 704602 110382 704838
rect 109826 704282 110062 704518
rect 110146 704282 110382 704518
rect 109826 687218 110062 687454
rect 110146 687218 110382 687454
rect 109826 686898 110062 687134
rect 110146 686898 110382 687134
rect 109826 651218 110062 651454
rect 110146 651218 110382 651454
rect 109826 650898 110062 651134
rect 110146 650898 110382 651134
rect 109826 615218 110062 615454
rect 110146 615218 110382 615454
rect 109826 614898 110062 615134
rect 110146 614898 110382 615134
rect 109826 579218 110062 579454
rect 110146 579218 110382 579454
rect 109826 578898 110062 579134
rect 110146 578898 110382 579134
rect 109826 543218 110062 543454
rect 110146 543218 110382 543454
rect 109826 542898 110062 543134
rect 110146 542898 110382 543134
rect 109826 507218 110062 507454
rect 110146 507218 110382 507454
rect 109826 506898 110062 507134
rect 110146 506898 110382 507134
rect 109826 471218 110062 471454
rect 110146 471218 110382 471454
rect 109826 470898 110062 471134
rect 110146 470898 110382 471134
rect 109826 435218 110062 435454
rect 110146 435218 110382 435454
rect 109826 434898 110062 435134
rect 110146 434898 110382 435134
rect 109826 399218 110062 399454
rect 110146 399218 110382 399454
rect 109826 398898 110062 399134
rect 110146 398898 110382 399134
rect 109826 363218 110062 363454
rect 110146 363218 110382 363454
rect 109826 362898 110062 363134
rect 110146 362898 110382 363134
rect 109826 327218 110062 327454
rect 110146 327218 110382 327454
rect 109826 326898 110062 327134
rect 110146 326898 110382 327134
rect 109826 291218 110062 291454
rect 110146 291218 110382 291454
rect 109826 290898 110062 291134
rect 110146 290898 110382 291134
rect 109826 255218 110062 255454
rect 110146 255218 110382 255454
rect 109826 254898 110062 255134
rect 110146 254898 110382 255134
rect 109826 219218 110062 219454
rect 110146 219218 110382 219454
rect 109826 218898 110062 219134
rect 110146 218898 110382 219134
rect 109826 183218 110062 183454
rect 110146 183218 110382 183454
rect 109826 182898 110062 183134
rect 110146 182898 110382 183134
rect 109826 147218 110062 147454
rect 110146 147218 110382 147454
rect 109826 146898 110062 147134
rect 110146 146898 110382 147134
rect 109826 111218 110062 111454
rect 110146 111218 110382 111454
rect 109826 110898 110062 111134
rect 110146 110898 110382 111134
rect 109826 75218 110062 75454
rect 110146 75218 110382 75454
rect 109826 74898 110062 75134
rect 110146 74898 110382 75134
rect 109826 39218 110062 39454
rect 110146 39218 110382 39454
rect 109826 38898 110062 39134
rect 110146 38898 110382 39134
rect 109826 3218 110062 3454
rect 110146 3218 110382 3454
rect 109826 2898 110062 3134
rect 110146 2898 110382 3134
rect 109826 -582 110062 -346
rect 110146 -582 110382 -346
rect 109826 -902 110062 -666
rect 110146 -902 110382 -666
rect 113546 690938 113782 691174
rect 113866 690938 114102 691174
rect 113546 690618 113782 690854
rect 113866 690618 114102 690854
rect 113546 654938 113782 655174
rect 113866 654938 114102 655174
rect 113546 654618 113782 654854
rect 113866 654618 114102 654854
rect 113546 618938 113782 619174
rect 113866 618938 114102 619174
rect 113546 618618 113782 618854
rect 113866 618618 114102 618854
rect 113546 582938 113782 583174
rect 113866 582938 114102 583174
rect 113546 582618 113782 582854
rect 113866 582618 114102 582854
rect 113546 546938 113782 547174
rect 113866 546938 114102 547174
rect 113546 546618 113782 546854
rect 113866 546618 114102 546854
rect 113546 510938 113782 511174
rect 113866 510938 114102 511174
rect 113546 510618 113782 510854
rect 113866 510618 114102 510854
rect 113546 474938 113782 475174
rect 113866 474938 114102 475174
rect 113546 474618 113782 474854
rect 113866 474618 114102 474854
rect 113546 438938 113782 439174
rect 113866 438938 114102 439174
rect 113546 438618 113782 438854
rect 113866 438618 114102 438854
rect 113546 402938 113782 403174
rect 113866 402938 114102 403174
rect 113546 402618 113782 402854
rect 113866 402618 114102 402854
rect 113546 366938 113782 367174
rect 113866 366938 114102 367174
rect 113546 366618 113782 366854
rect 113866 366618 114102 366854
rect 113546 330938 113782 331174
rect 113866 330938 114102 331174
rect 113546 330618 113782 330854
rect 113866 330618 114102 330854
rect 113546 294938 113782 295174
rect 113866 294938 114102 295174
rect 113546 294618 113782 294854
rect 113866 294618 114102 294854
rect 113546 258938 113782 259174
rect 113866 258938 114102 259174
rect 113546 258618 113782 258854
rect 113866 258618 114102 258854
rect 113546 222938 113782 223174
rect 113866 222938 114102 223174
rect 113546 222618 113782 222854
rect 113866 222618 114102 222854
rect 113546 186938 113782 187174
rect 113866 186938 114102 187174
rect 113546 186618 113782 186854
rect 113866 186618 114102 186854
rect 113546 150938 113782 151174
rect 113866 150938 114102 151174
rect 113546 150618 113782 150854
rect 113866 150618 114102 150854
rect 113546 114938 113782 115174
rect 113866 114938 114102 115174
rect 113546 114618 113782 114854
rect 113866 114618 114102 114854
rect 113546 78938 113782 79174
rect 113866 78938 114102 79174
rect 113546 78618 113782 78854
rect 113866 78618 114102 78854
rect 113546 42938 113782 43174
rect 113866 42938 114102 43174
rect 113546 42618 113782 42854
rect 113866 42618 114102 42854
rect 113546 6938 113782 7174
rect 113866 6938 114102 7174
rect 113546 6618 113782 6854
rect 113866 6618 114102 6854
rect 113546 -2502 113782 -2266
rect 113866 -2502 114102 -2266
rect 113546 -2822 113782 -2586
rect 113866 -2822 114102 -2586
rect 117266 694658 117502 694894
rect 117586 694658 117822 694894
rect 117266 694338 117502 694574
rect 117586 694338 117822 694574
rect 117266 658658 117502 658894
rect 117586 658658 117822 658894
rect 117266 658338 117502 658574
rect 117586 658338 117822 658574
rect 117266 622658 117502 622894
rect 117586 622658 117822 622894
rect 117266 622338 117502 622574
rect 117586 622338 117822 622574
rect 117266 586658 117502 586894
rect 117586 586658 117822 586894
rect 117266 586338 117502 586574
rect 117586 586338 117822 586574
rect 117266 550658 117502 550894
rect 117586 550658 117822 550894
rect 117266 550338 117502 550574
rect 117586 550338 117822 550574
rect 117266 514658 117502 514894
rect 117586 514658 117822 514894
rect 117266 514338 117502 514574
rect 117586 514338 117822 514574
rect 117266 478658 117502 478894
rect 117586 478658 117822 478894
rect 117266 478338 117502 478574
rect 117586 478338 117822 478574
rect 117266 442658 117502 442894
rect 117586 442658 117822 442894
rect 117266 442338 117502 442574
rect 117586 442338 117822 442574
rect 117266 406658 117502 406894
rect 117586 406658 117822 406894
rect 117266 406338 117502 406574
rect 117586 406338 117822 406574
rect 117266 370658 117502 370894
rect 117586 370658 117822 370894
rect 117266 370338 117502 370574
rect 117586 370338 117822 370574
rect 117266 334658 117502 334894
rect 117586 334658 117822 334894
rect 117266 334338 117502 334574
rect 117586 334338 117822 334574
rect 117266 298658 117502 298894
rect 117586 298658 117822 298894
rect 117266 298338 117502 298574
rect 117586 298338 117822 298574
rect 117266 262658 117502 262894
rect 117586 262658 117822 262894
rect 117266 262338 117502 262574
rect 117586 262338 117822 262574
rect 117266 226658 117502 226894
rect 117586 226658 117822 226894
rect 117266 226338 117502 226574
rect 117586 226338 117822 226574
rect 117266 190658 117502 190894
rect 117586 190658 117822 190894
rect 117266 190338 117502 190574
rect 117586 190338 117822 190574
rect 117266 154658 117502 154894
rect 117586 154658 117822 154894
rect 117266 154338 117502 154574
rect 117586 154338 117822 154574
rect 117266 118658 117502 118894
rect 117586 118658 117822 118894
rect 117266 118338 117502 118574
rect 117586 118338 117822 118574
rect 117266 82658 117502 82894
rect 117586 82658 117822 82894
rect 117266 82338 117502 82574
rect 117586 82338 117822 82574
rect 117266 46658 117502 46894
rect 117586 46658 117822 46894
rect 117266 46338 117502 46574
rect 117586 46338 117822 46574
rect 117266 10658 117502 10894
rect 117586 10658 117822 10894
rect 117266 10338 117502 10574
rect 117586 10338 117822 10574
rect 117266 -4422 117502 -4186
rect 117586 -4422 117822 -4186
rect 117266 -4742 117502 -4506
rect 117586 -4742 117822 -4506
rect 138986 711322 139222 711558
rect 139306 711322 139542 711558
rect 138986 711002 139222 711238
rect 139306 711002 139542 711238
rect 135266 709402 135502 709638
rect 135586 709402 135822 709638
rect 135266 709082 135502 709318
rect 135586 709082 135822 709318
rect 131546 707482 131782 707718
rect 131866 707482 132102 707718
rect 131546 707162 131782 707398
rect 131866 707162 132102 707398
rect 120986 698378 121222 698614
rect 121306 698378 121542 698614
rect 120986 698058 121222 698294
rect 121306 698058 121542 698294
rect 120986 662378 121222 662614
rect 121306 662378 121542 662614
rect 120986 662058 121222 662294
rect 121306 662058 121542 662294
rect 120986 626378 121222 626614
rect 121306 626378 121542 626614
rect 120986 626058 121222 626294
rect 121306 626058 121542 626294
rect 120986 590378 121222 590614
rect 121306 590378 121542 590614
rect 120986 590058 121222 590294
rect 121306 590058 121542 590294
rect 120986 554378 121222 554614
rect 121306 554378 121542 554614
rect 120986 554058 121222 554294
rect 121306 554058 121542 554294
rect 120986 518378 121222 518614
rect 121306 518378 121542 518614
rect 120986 518058 121222 518294
rect 121306 518058 121542 518294
rect 120986 482378 121222 482614
rect 121306 482378 121542 482614
rect 120986 482058 121222 482294
rect 121306 482058 121542 482294
rect 120986 446378 121222 446614
rect 121306 446378 121542 446614
rect 120986 446058 121222 446294
rect 121306 446058 121542 446294
rect 120986 410378 121222 410614
rect 121306 410378 121542 410614
rect 120986 410058 121222 410294
rect 121306 410058 121542 410294
rect 120986 374378 121222 374614
rect 121306 374378 121542 374614
rect 120986 374058 121222 374294
rect 121306 374058 121542 374294
rect 120986 338378 121222 338614
rect 121306 338378 121542 338614
rect 120986 338058 121222 338294
rect 121306 338058 121542 338294
rect 120986 302378 121222 302614
rect 121306 302378 121542 302614
rect 120986 302058 121222 302294
rect 121306 302058 121542 302294
rect 120986 266378 121222 266614
rect 121306 266378 121542 266614
rect 120986 266058 121222 266294
rect 121306 266058 121542 266294
rect 120986 230378 121222 230614
rect 121306 230378 121542 230614
rect 120986 230058 121222 230294
rect 121306 230058 121542 230294
rect 120986 194378 121222 194614
rect 121306 194378 121542 194614
rect 120986 194058 121222 194294
rect 121306 194058 121542 194294
rect 120986 158378 121222 158614
rect 121306 158378 121542 158614
rect 120986 158058 121222 158294
rect 121306 158058 121542 158294
rect 120986 122378 121222 122614
rect 121306 122378 121542 122614
rect 120986 122058 121222 122294
rect 121306 122058 121542 122294
rect 120986 86378 121222 86614
rect 121306 86378 121542 86614
rect 120986 86058 121222 86294
rect 121306 86058 121542 86294
rect 120986 50378 121222 50614
rect 121306 50378 121542 50614
rect 120986 50058 121222 50294
rect 121306 50058 121542 50294
rect 120986 14378 121222 14614
rect 121306 14378 121542 14614
rect 120986 14058 121222 14294
rect 121306 14058 121542 14294
rect 102986 -7302 103222 -7066
rect 103306 -7302 103542 -7066
rect 102986 -7622 103222 -7386
rect 103306 -7622 103542 -7386
rect 127826 705562 128062 705798
rect 128146 705562 128382 705798
rect 127826 705242 128062 705478
rect 128146 705242 128382 705478
rect 127826 669218 128062 669454
rect 128146 669218 128382 669454
rect 127826 668898 128062 669134
rect 128146 668898 128382 669134
rect 127826 633218 128062 633454
rect 128146 633218 128382 633454
rect 127826 632898 128062 633134
rect 128146 632898 128382 633134
rect 127826 597218 128062 597454
rect 128146 597218 128382 597454
rect 127826 596898 128062 597134
rect 128146 596898 128382 597134
rect 127826 561218 128062 561454
rect 128146 561218 128382 561454
rect 127826 560898 128062 561134
rect 128146 560898 128382 561134
rect 127826 525218 128062 525454
rect 128146 525218 128382 525454
rect 127826 524898 128062 525134
rect 128146 524898 128382 525134
rect 127826 489218 128062 489454
rect 128146 489218 128382 489454
rect 127826 488898 128062 489134
rect 128146 488898 128382 489134
rect 127826 453218 128062 453454
rect 128146 453218 128382 453454
rect 127826 452898 128062 453134
rect 128146 452898 128382 453134
rect 127826 417218 128062 417454
rect 128146 417218 128382 417454
rect 127826 416898 128062 417134
rect 128146 416898 128382 417134
rect 127826 381218 128062 381454
rect 128146 381218 128382 381454
rect 127826 380898 128062 381134
rect 128146 380898 128382 381134
rect 127826 345218 128062 345454
rect 128146 345218 128382 345454
rect 127826 344898 128062 345134
rect 128146 344898 128382 345134
rect 127826 309218 128062 309454
rect 128146 309218 128382 309454
rect 127826 308898 128062 309134
rect 128146 308898 128382 309134
rect 127826 273218 128062 273454
rect 128146 273218 128382 273454
rect 127826 272898 128062 273134
rect 128146 272898 128382 273134
rect 127826 237218 128062 237454
rect 128146 237218 128382 237454
rect 127826 236898 128062 237134
rect 128146 236898 128382 237134
rect 127826 201218 128062 201454
rect 128146 201218 128382 201454
rect 127826 200898 128062 201134
rect 128146 200898 128382 201134
rect 127826 165218 128062 165454
rect 128146 165218 128382 165454
rect 127826 164898 128062 165134
rect 128146 164898 128382 165134
rect 127826 129218 128062 129454
rect 128146 129218 128382 129454
rect 127826 128898 128062 129134
rect 128146 128898 128382 129134
rect 127826 93218 128062 93454
rect 128146 93218 128382 93454
rect 127826 92898 128062 93134
rect 128146 92898 128382 93134
rect 127826 57218 128062 57454
rect 128146 57218 128382 57454
rect 127826 56898 128062 57134
rect 128146 56898 128382 57134
rect 127826 21218 128062 21454
rect 128146 21218 128382 21454
rect 127826 20898 128062 21134
rect 128146 20898 128382 21134
rect 127826 -1542 128062 -1306
rect 128146 -1542 128382 -1306
rect 127826 -1862 128062 -1626
rect 128146 -1862 128382 -1626
rect 131546 672938 131782 673174
rect 131866 672938 132102 673174
rect 131546 672618 131782 672854
rect 131866 672618 132102 672854
rect 131546 636938 131782 637174
rect 131866 636938 132102 637174
rect 131546 636618 131782 636854
rect 131866 636618 132102 636854
rect 131546 600938 131782 601174
rect 131866 600938 132102 601174
rect 131546 600618 131782 600854
rect 131866 600618 132102 600854
rect 131546 564938 131782 565174
rect 131866 564938 132102 565174
rect 131546 564618 131782 564854
rect 131866 564618 132102 564854
rect 131546 528938 131782 529174
rect 131866 528938 132102 529174
rect 131546 528618 131782 528854
rect 131866 528618 132102 528854
rect 131546 492938 131782 493174
rect 131866 492938 132102 493174
rect 131546 492618 131782 492854
rect 131866 492618 132102 492854
rect 131546 456938 131782 457174
rect 131866 456938 132102 457174
rect 131546 456618 131782 456854
rect 131866 456618 132102 456854
rect 131546 420938 131782 421174
rect 131866 420938 132102 421174
rect 131546 420618 131782 420854
rect 131866 420618 132102 420854
rect 131546 384938 131782 385174
rect 131866 384938 132102 385174
rect 131546 384618 131782 384854
rect 131866 384618 132102 384854
rect 131546 348938 131782 349174
rect 131866 348938 132102 349174
rect 131546 348618 131782 348854
rect 131866 348618 132102 348854
rect 131546 312938 131782 313174
rect 131866 312938 132102 313174
rect 131546 312618 131782 312854
rect 131866 312618 132102 312854
rect 131546 276938 131782 277174
rect 131866 276938 132102 277174
rect 131546 276618 131782 276854
rect 131866 276618 132102 276854
rect 131546 240938 131782 241174
rect 131866 240938 132102 241174
rect 131546 240618 131782 240854
rect 131866 240618 132102 240854
rect 131546 204938 131782 205174
rect 131866 204938 132102 205174
rect 131546 204618 131782 204854
rect 131866 204618 132102 204854
rect 131546 168938 131782 169174
rect 131866 168938 132102 169174
rect 131546 168618 131782 168854
rect 131866 168618 132102 168854
rect 131546 132938 131782 133174
rect 131866 132938 132102 133174
rect 131546 132618 131782 132854
rect 131866 132618 132102 132854
rect 131546 96938 131782 97174
rect 131866 96938 132102 97174
rect 131546 96618 131782 96854
rect 131866 96618 132102 96854
rect 131546 60938 131782 61174
rect 131866 60938 132102 61174
rect 131546 60618 131782 60854
rect 131866 60618 132102 60854
rect 131546 24938 131782 25174
rect 131866 24938 132102 25174
rect 131546 24618 131782 24854
rect 131866 24618 132102 24854
rect 131546 -3462 131782 -3226
rect 131866 -3462 132102 -3226
rect 131546 -3782 131782 -3546
rect 131866 -3782 132102 -3546
rect 135266 676658 135502 676894
rect 135586 676658 135822 676894
rect 135266 676338 135502 676574
rect 135586 676338 135822 676574
rect 135266 640658 135502 640894
rect 135586 640658 135822 640894
rect 135266 640338 135502 640574
rect 135586 640338 135822 640574
rect 135266 604658 135502 604894
rect 135586 604658 135822 604894
rect 135266 604338 135502 604574
rect 135586 604338 135822 604574
rect 135266 568658 135502 568894
rect 135586 568658 135822 568894
rect 135266 568338 135502 568574
rect 135586 568338 135822 568574
rect 135266 532658 135502 532894
rect 135586 532658 135822 532894
rect 135266 532338 135502 532574
rect 135586 532338 135822 532574
rect 135266 496658 135502 496894
rect 135586 496658 135822 496894
rect 135266 496338 135502 496574
rect 135586 496338 135822 496574
rect 135266 460658 135502 460894
rect 135586 460658 135822 460894
rect 135266 460338 135502 460574
rect 135586 460338 135822 460574
rect 135266 424658 135502 424894
rect 135586 424658 135822 424894
rect 135266 424338 135502 424574
rect 135586 424338 135822 424574
rect 135266 388658 135502 388894
rect 135586 388658 135822 388894
rect 135266 388338 135502 388574
rect 135586 388338 135822 388574
rect 135266 352658 135502 352894
rect 135586 352658 135822 352894
rect 135266 352338 135502 352574
rect 135586 352338 135822 352574
rect 135266 316658 135502 316894
rect 135586 316658 135822 316894
rect 135266 316338 135502 316574
rect 135586 316338 135822 316574
rect 135266 280658 135502 280894
rect 135586 280658 135822 280894
rect 135266 280338 135502 280574
rect 135586 280338 135822 280574
rect 135266 244658 135502 244894
rect 135586 244658 135822 244894
rect 135266 244338 135502 244574
rect 135586 244338 135822 244574
rect 135266 208658 135502 208894
rect 135586 208658 135822 208894
rect 135266 208338 135502 208574
rect 135586 208338 135822 208574
rect 135266 172658 135502 172894
rect 135586 172658 135822 172894
rect 135266 172338 135502 172574
rect 135586 172338 135822 172574
rect 135266 136658 135502 136894
rect 135586 136658 135822 136894
rect 135266 136338 135502 136574
rect 135586 136338 135822 136574
rect 135266 100658 135502 100894
rect 135586 100658 135822 100894
rect 135266 100338 135502 100574
rect 135586 100338 135822 100574
rect 135266 64658 135502 64894
rect 135586 64658 135822 64894
rect 135266 64338 135502 64574
rect 135586 64338 135822 64574
rect 135266 28658 135502 28894
rect 135586 28658 135822 28894
rect 135266 28338 135502 28574
rect 135586 28338 135822 28574
rect 135266 -5382 135502 -5146
rect 135586 -5382 135822 -5146
rect 135266 -5702 135502 -5466
rect 135586 -5702 135822 -5466
rect 156986 710362 157222 710598
rect 157306 710362 157542 710598
rect 156986 710042 157222 710278
rect 157306 710042 157542 710278
rect 153266 708442 153502 708678
rect 153586 708442 153822 708678
rect 153266 708122 153502 708358
rect 153586 708122 153822 708358
rect 149546 706522 149782 706758
rect 149866 706522 150102 706758
rect 149546 706202 149782 706438
rect 149866 706202 150102 706438
rect 138986 680378 139222 680614
rect 139306 680378 139542 680614
rect 138986 680058 139222 680294
rect 139306 680058 139542 680294
rect 138986 644378 139222 644614
rect 139306 644378 139542 644614
rect 138986 644058 139222 644294
rect 139306 644058 139542 644294
rect 138986 608378 139222 608614
rect 139306 608378 139542 608614
rect 138986 608058 139222 608294
rect 139306 608058 139542 608294
rect 138986 572378 139222 572614
rect 139306 572378 139542 572614
rect 138986 572058 139222 572294
rect 139306 572058 139542 572294
rect 138986 536378 139222 536614
rect 139306 536378 139542 536614
rect 138986 536058 139222 536294
rect 139306 536058 139542 536294
rect 138986 500378 139222 500614
rect 139306 500378 139542 500614
rect 138986 500058 139222 500294
rect 139306 500058 139542 500294
rect 138986 464378 139222 464614
rect 139306 464378 139542 464614
rect 138986 464058 139222 464294
rect 139306 464058 139542 464294
rect 138986 428378 139222 428614
rect 139306 428378 139542 428614
rect 138986 428058 139222 428294
rect 139306 428058 139542 428294
rect 138986 392378 139222 392614
rect 139306 392378 139542 392614
rect 138986 392058 139222 392294
rect 139306 392058 139542 392294
rect 138986 356378 139222 356614
rect 139306 356378 139542 356614
rect 138986 356058 139222 356294
rect 139306 356058 139542 356294
rect 138986 320378 139222 320614
rect 139306 320378 139542 320614
rect 138986 320058 139222 320294
rect 139306 320058 139542 320294
rect 138986 284378 139222 284614
rect 139306 284378 139542 284614
rect 138986 284058 139222 284294
rect 139306 284058 139542 284294
rect 138986 248378 139222 248614
rect 139306 248378 139542 248614
rect 138986 248058 139222 248294
rect 139306 248058 139542 248294
rect 138986 212378 139222 212614
rect 139306 212378 139542 212614
rect 138986 212058 139222 212294
rect 139306 212058 139542 212294
rect 138986 176378 139222 176614
rect 139306 176378 139542 176614
rect 138986 176058 139222 176294
rect 139306 176058 139542 176294
rect 138986 140378 139222 140614
rect 139306 140378 139542 140614
rect 138986 140058 139222 140294
rect 139306 140058 139542 140294
rect 138986 104378 139222 104614
rect 139306 104378 139542 104614
rect 138986 104058 139222 104294
rect 139306 104058 139542 104294
rect 138986 68378 139222 68614
rect 139306 68378 139542 68614
rect 138986 68058 139222 68294
rect 139306 68058 139542 68294
rect 138986 32378 139222 32614
rect 139306 32378 139542 32614
rect 138986 32058 139222 32294
rect 139306 32058 139542 32294
rect 120986 -6342 121222 -6106
rect 121306 -6342 121542 -6106
rect 120986 -6662 121222 -6426
rect 121306 -6662 121542 -6426
rect 145826 704602 146062 704838
rect 146146 704602 146382 704838
rect 145826 704282 146062 704518
rect 146146 704282 146382 704518
rect 145826 687218 146062 687454
rect 146146 687218 146382 687454
rect 145826 686898 146062 687134
rect 146146 686898 146382 687134
rect 145826 651218 146062 651454
rect 146146 651218 146382 651454
rect 145826 650898 146062 651134
rect 146146 650898 146382 651134
rect 145826 615218 146062 615454
rect 146146 615218 146382 615454
rect 145826 614898 146062 615134
rect 146146 614898 146382 615134
rect 145826 579218 146062 579454
rect 146146 579218 146382 579454
rect 145826 578898 146062 579134
rect 146146 578898 146382 579134
rect 145826 543218 146062 543454
rect 146146 543218 146382 543454
rect 145826 542898 146062 543134
rect 146146 542898 146382 543134
rect 145826 507218 146062 507454
rect 146146 507218 146382 507454
rect 145826 506898 146062 507134
rect 146146 506898 146382 507134
rect 145826 471218 146062 471454
rect 146146 471218 146382 471454
rect 145826 470898 146062 471134
rect 146146 470898 146382 471134
rect 145826 435218 146062 435454
rect 146146 435218 146382 435454
rect 145826 434898 146062 435134
rect 146146 434898 146382 435134
rect 145826 399218 146062 399454
rect 146146 399218 146382 399454
rect 145826 398898 146062 399134
rect 146146 398898 146382 399134
rect 145826 363218 146062 363454
rect 146146 363218 146382 363454
rect 145826 362898 146062 363134
rect 146146 362898 146382 363134
rect 145826 327218 146062 327454
rect 146146 327218 146382 327454
rect 145826 326898 146062 327134
rect 146146 326898 146382 327134
rect 145826 291218 146062 291454
rect 146146 291218 146382 291454
rect 145826 290898 146062 291134
rect 146146 290898 146382 291134
rect 145826 255218 146062 255454
rect 146146 255218 146382 255454
rect 145826 254898 146062 255134
rect 146146 254898 146382 255134
rect 145826 219218 146062 219454
rect 146146 219218 146382 219454
rect 145826 218898 146062 219134
rect 146146 218898 146382 219134
rect 145826 183218 146062 183454
rect 146146 183218 146382 183454
rect 145826 182898 146062 183134
rect 146146 182898 146382 183134
rect 145826 147218 146062 147454
rect 146146 147218 146382 147454
rect 145826 146898 146062 147134
rect 146146 146898 146382 147134
rect 145826 111218 146062 111454
rect 146146 111218 146382 111454
rect 145826 110898 146062 111134
rect 146146 110898 146382 111134
rect 145826 75218 146062 75454
rect 146146 75218 146382 75454
rect 145826 74898 146062 75134
rect 146146 74898 146382 75134
rect 145826 39218 146062 39454
rect 146146 39218 146382 39454
rect 145826 38898 146062 39134
rect 146146 38898 146382 39134
rect 145826 3218 146062 3454
rect 146146 3218 146382 3454
rect 145826 2898 146062 3134
rect 146146 2898 146382 3134
rect 145826 -582 146062 -346
rect 146146 -582 146382 -346
rect 145826 -902 146062 -666
rect 146146 -902 146382 -666
rect 149546 690938 149782 691174
rect 149866 690938 150102 691174
rect 149546 690618 149782 690854
rect 149866 690618 150102 690854
rect 149546 654938 149782 655174
rect 149866 654938 150102 655174
rect 149546 654618 149782 654854
rect 149866 654618 150102 654854
rect 149546 618938 149782 619174
rect 149866 618938 150102 619174
rect 149546 618618 149782 618854
rect 149866 618618 150102 618854
rect 149546 582938 149782 583174
rect 149866 582938 150102 583174
rect 149546 582618 149782 582854
rect 149866 582618 150102 582854
rect 149546 546938 149782 547174
rect 149866 546938 150102 547174
rect 149546 546618 149782 546854
rect 149866 546618 150102 546854
rect 149546 510938 149782 511174
rect 149866 510938 150102 511174
rect 149546 510618 149782 510854
rect 149866 510618 150102 510854
rect 149546 474938 149782 475174
rect 149866 474938 150102 475174
rect 149546 474618 149782 474854
rect 149866 474618 150102 474854
rect 149546 438938 149782 439174
rect 149866 438938 150102 439174
rect 149546 438618 149782 438854
rect 149866 438618 150102 438854
rect 149546 402938 149782 403174
rect 149866 402938 150102 403174
rect 149546 402618 149782 402854
rect 149866 402618 150102 402854
rect 149546 366938 149782 367174
rect 149866 366938 150102 367174
rect 149546 366618 149782 366854
rect 149866 366618 150102 366854
rect 149546 330938 149782 331174
rect 149866 330938 150102 331174
rect 149546 330618 149782 330854
rect 149866 330618 150102 330854
rect 149546 294938 149782 295174
rect 149866 294938 150102 295174
rect 149546 294618 149782 294854
rect 149866 294618 150102 294854
rect 149546 258938 149782 259174
rect 149866 258938 150102 259174
rect 149546 258618 149782 258854
rect 149866 258618 150102 258854
rect 149546 222938 149782 223174
rect 149866 222938 150102 223174
rect 149546 222618 149782 222854
rect 149866 222618 150102 222854
rect 149546 186938 149782 187174
rect 149866 186938 150102 187174
rect 149546 186618 149782 186854
rect 149866 186618 150102 186854
rect 149546 150938 149782 151174
rect 149866 150938 150102 151174
rect 149546 150618 149782 150854
rect 149866 150618 150102 150854
rect 149546 114938 149782 115174
rect 149866 114938 150102 115174
rect 149546 114618 149782 114854
rect 149866 114618 150102 114854
rect 149546 78938 149782 79174
rect 149866 78938 150102 79174
rect 149546 78618 149782 78854
rect 149866 78618 150102 78854
rect 149546 42938 149782 43174
rect 149866 42938 150102 43174
rect 149546 42618 149782 42854
rect 149866 42618 150102 42854
rect 149546 6938 149782 7174
rect 149866 6938 150102 7174
rect 149546 6618 149782 6854
rect 149866 6618 150102 6854
rect 149546 -2502 149782 -2266
rect 149866 -2502 150102 -2266
rect 149546 -2822 149782 -2586
rect 149866 -2822 150102 -2586
rect 153266 694658 153502 694894
rect 153586 694658 153822 694894
rect 153266 694338 153502 694574
rect 153586 694338 153822 694574
rect 153266 658658 153502 658894
rect 153586 658658 153822 658894
rect 153266 658338 153502 658574
rect 153586 658338 153822 658574
rect 153266 622658 153502 622894
rect 153586 622658 153822 622894
rect 153266 622338 153502 622574
rect 153586 622338 153822 622574
rect 153266 586658 153502 586894
rect 153586 586658 153822 586894
rect 153266 586338 153502 586574
rect 153586 586338 153822 586574
rect 153266 550658 153502 550894
rect 153586 550658 153822 550894
rect 153266 550338 153502 550574
rect 153586 550338 153822 550574
rect 153266 514658 153502 514894
rect 153586 514658 153822 514894
rect 153266 514338 153502 514574
rect 153586 514338 153822 514574
rect 153266 478658 153502 478894
rect 153586 478658 153822 478894
rect 153266 478338 153502 478574
rect 153586 478338 153822 478574
rect 153266 442658 153502 442894
rect 153586 442658 153822 442894
rect 153266 442338 153502 442574
rect 153586 442338 153822 442574
rect 153266 406658 153502 406894
rect 153586 406658 153822 406894
rect 153266 406338 153502 406574
rect 153586 406338 153822 406574
rect 153266 370658 153502 370894
rect 153586 370658 153822 370894
rect 153266 370338 153502 370574
rect 153586 370338 153822 370574
rect 153266 334658 153502 334894
rect 153586 334658 153822 334894
rect 153266 334338 153502 334574
rect 153586 334338 153822 334574
rect 153266 298658 153502 298894
rect 153586 298658 153822 298894
rect 153266 298338 153502 298574
rect 153586 298338 153822 298574
rect 153266 262658 153502 262894
rect 153586 262658 153822 262894
rect 153266 262338 153502 262574
rect 153586 262338 153822 262574
rect 153266 226658 153502 226894
rect 153586 226658 153822 226894
rect 153266 226338 153502 226574
rect 153586 226338 153822 226574
rect 153266 190658 153502 190894
rect 153586 190658 153822 190894
rect 153266 190338 153502 190574
rect 153586 190338 153822 190574
rect 153266 154658 153502 154894
rect 153586 154658 153822 154894
rect 153266 154338 153502 154574
rect 153586 154338 153822 154574
rect 153266 118658 153502 118894
rect 153586 118658 153822 118894
rect 153266 118338 153502 118574
rect 153586 118338 153822 118574
rect 153266 82658 153502 82894
rect 153586 82658 153822 82894
rect 153266 82338 153502 82574
rect 153586 82338 153822 82574
rect 153266 46658 153502 46894
rect 153586 46658 153822 46894
rect 153266 46338 153502 46574
rect 153586 46338 153822 46574
rect 153266 10658 153502 10894
rect 153586 10658 153822 10894
rect 153266 10338 153502 10574
rect 153586 10338 153822 10574
rect 153266 -4422 153502 -4186
rect 153586 -4422 153822 -4186
rect 153266 -4742 153502 -4506
rect 153586 -4742 153822 -4506
rect 174986 711322 175222 711558
rect 175306 711322 175542 711558
rect 174986 711002 175222 711238
rect 175306 711002 175542 711238
rect 171266 709402 171502 709638
rect 171586 709402 171822 709638
rect 171266 709082 171502 709318
rect 171586 709082 171822 709318
rect 167546 707482 167782 707718
rect 167866 707482 168102 707718
rect 167546 707162 167782 707398
rect 167866 707162 168102 707398
rect 156986 698378 157222 698614
rect 157306 698378 157542 698614
rect 156986 698058 157222 698294
rect 157306 698058 157542 698294
rect 156986 662378 157222 662614
rect 157306 662378 157542 662614
rect 156986 662058 157222 662294
rect 157306 662058 157542 662294
rect 156986 626378 157222 626614
rect 157306 626378 157542 626614
rect 156986 626058 157222 626294
rect 157306 626058 157542 626294
rect 156986 590378 157222 590614
rect 157306 590378 157542 590614
rect 156986 590058 157222 590294
rect 157306 590058 157542 590294
rect 156986 554378 157222 554614
rect 157306 554378 157542 554614
rect 156986 554058 157222 554294
rect 157306 554058 157542 554294
rect 156986 518378 157222 518614
rect 157306 518378 157542 518614
rect 156986 518058 157222 518294
rect 157306 518058 157542 518294
rect 163826 705562 164062 705798
rect 164146 705562 164382 705798
rect 163826 705242 164062 705478
rect 164146 705242 164382 705478
rect 163826 669218 164062 669454
rect 164146 669218 164382 669454
rect 163826 668898 164062 669134
rect 164146 668898 164382 669134
rect 163826 633218 164062 633454
rect 164146 633218 164382 633454
rect 163826 632898 164062 633134
rect 164146 632898 164382 633134
rect 163826 597218 164062 597454
rect 164146 597218 164382 597454
rect 163826 596898 164062 597134
rect 164146 596898 164382 597134
rect 163826 561218 164062 561454
rect 164146 561218 164382 561454
rect 163826 560898 164062 561134
rect 164146 560898 164382 561134
rect 163826 525218 164062 525454
rect 164146 525218 164382 525454
rect 163826 524898 164062 525134
rect 164146 524898 164382 525134
rect 167546 672938 167782 673174
rect 167866 672938 168102 673174
rect 167546 672618 167782 672854
rect 167866 672618 168102 672854
rect 167546 636938 167782 637174
rect 167866 636938 168102 637174
rect 167546 636618 167782 636854
rect 167866 636618 168102 636854
rect 167546 600938 167782 601174
rect 167866 600938 168102 601174
rect 167546 600618 167782 600854
rect 167866 600618 168102 600854
rect 167546 564938 167782 565174
rect 167866 564938 168102 565174
rect 167546 564618 167782 564854
rect 167866 564618 168102 564854
rect 167546 528938 167782 529174
rect 167866 528938 168102 529174
rect 167546 528618 167782 528854
rect 167866 528618 168102 528854
rect 171266 676658 171502 676894
rect 171586 676658 171822 676894
rect 171266 676338 171502 676574
rect 171586 676338 171822 676574
rect 171266 640658 171502 640894
rect 171586 640658 171822 640894
rect 171266 640338 171502 640574
rect 171586 640338 171822 640574
rect 171266 604658 171502 604894
rect 171586 604658 171822 604894
rect 171266 604338 171502 604574
rect 171586 604338 171822 604574
rect 171266 568658 171502 568894
rect 171586 568658 171822 568894
rect 171266 568338 171502 568574
rect 171586 568338 171822 568574
rect 171266 532658 171502 532894
rect 171586 532658 171822 532894
rect 171266 532338 171502 532574
rect 171586 532338 171822 532574
rect 192986 710362 193222 710598
rect 193306 710362 193542 710598
rect 192986 710042 193222 710278
rect 193306 710042 193542 710278
rect 189266 708442 189502 708678
rect 189586 708442 189822 708678
rect 189266 708122 189502 708358
rect 189586 708122 189822 708358
rect 185546 706522 185782 706758
rect 185866 706522 186102 706758
rect 185546 706202 185782 706438
rect 185866 706202 186102 706438
rect 174986 680378 175222 680614
rect 175306 680378 175542 680614
rect 174986 680058 175222 680294
rect 175306 680058 175542 680294
rect 174986 644378 175222 644614
rect 175306 644378 175542 644614
rect 174986 644058 175222 644294
rect 175306 644058 175542 644294
rect 174986 608378 175222 608614
rect 175306 608378 175542 608614
rect 174986 608058 175222 608294
rect 175306 608058 175542 608294
rect 174986 572378 175222 572614
rect 175306 572378 175542 572614
rect 174986 572058 175222 572294
rect 175306 572058 175542 572294
rect 174986 536378 175222 536614
rect 175306 536378 175542 536614
rect 174986 536058 175222 536294
rect 175306 536058 175542 536294
rect 181826 704602 182062 704838
rect 182146 704602 182382 704838
rect 181826 704282 182062 704518
rect 182146 704282 182382 704518
rect 181826 687218 182062 687454
rect 182146 687218 182382 687454
rect 181826 686898 182062 687134
rect 182146 686898 182382 687134
rect 181826 651218 182062 651454
rect 182146 651218 182382 651454
rect 181826 650898 182062 651134
rect 182146 650898 182382 651134
rect 181826 615218 182062 615454
rect 182146 615218 182382 615454
rect 181826 614898 182062 615134
rect 182146 614898 182382 615134
rect 181826 579218 182062 579454
rect 182146 579218 182382 579454
rect 181826 578898 182062 579134
rect 182146 578898 182382 579134
rect 181826 543218 182062 543454
rect 182146 543218 182382 543454
rect 181826 542898 182062 543134
rect 182146 542898 182382 543134
rect 185546 690938 185782 691174
rect 185866 690938 186102 691174
rect 185546 690618 185782 690854
rect 185866 690618 186102 690854
rect 185546 654938 185782 655174
rect 185866 654938 186102 655174
rect 185546 654618 185782 654854
rect 185866 654618 186102 654854
rect 185546 618938 185782 619174
rect 185866 618938 186102 619174
rect 185546 618618 185782 618854
rect 185866 618618 186102 618854
rect 185546 582938 185782 583174
rect 185866 582938 186102 583174
rect 185546 582618 185782 582854
rect 185866 582618 186102 582854
rect 185546 546938 185782 547174
rect 185866 546938 186102 547174
rect 185546 546618 185782 546854
rect 185866 546618 186102 546854
rect 185546 510938 185782 511174
rect 185866 510938 186102 511174
rect 185546 510618 185782 510854
rect 185866 510618 186102 510854
rect 189266 694658 189502 694894
rect 189586 694658 189822 694894
rect 189266 694338 189502 694574
rect 189586 694338 189822 694574
rect 189266 658658 189502 658894
rect 189586 658658 189822 658894
rect 189266 658338 189502 658574
rect 189586 658338 189822 658574
rect 189266 622658 189502 622894
rect 189586 622658 189822 622894
rect 189266 622338 189502 622574
rect 189586 622338 189822 622574
rect 189266 586658 189502 586894
rect 189586 586658 189822 586894
rect 189266 586338 189502 586574
rect 189586 586338 189822 586574
rect 189266 550658 189502 550894
rect 189586 550658 189822 550894
rect 189266 550338 189502 550574
rect 189586 550338 189822 550574
rect 189266 514658 189502 514894
rect 189586 514658 189822 514894
rect 189266 514338 189502 514574
rect 189586 514338 189822 514574
rect 210986 711322 211222 711558
rect 211306 711322 211542 711558
rect 210986 711002 211222 711238
rect 211306 711002 211542 711238
rect 207266 709402 207502 709638
rect 207586 709402 207822 709638
rect 207266 709082 207502 709318
rect 207586 709082 207822 709318
rect 203546 707482 203782 707718
rect 203866 707482 204102 707718
rect 203546 707162 203782 707398
rect 203866 707162 204102 707398
rect 192986 698378 193222 698614
rect 193306 698378 193542 698614
rect 192986 698058 193222 698294
rect 193306 698058 193542 698294
rect 192986 662378 193222 662614
rect 193306 662378 193542 662614
rect 192986 662058 193222 662294
rect 193306 662058 193542 662294
rect 192986 626378 193222 626614
rect 193306 626378 193542 626614
rect 192986 626058 193222 626294
rect 193306 626058 193542 626294
rect 192986 590378 193222 590614
rect 193306 590378 193542 590614
rect 192986 590058 193222 590294
rect 193306 590058 193542 590294
rect 192986 554378 193222 554614
rect 193306 554378 193542 554614
rect 192986 554058 193222 554294
rect 193306 554058 193542 554294
rect 192986 518378 193222 518614
rect 193306 518378 193542 518614
rect 192986 518058 193222 518294
rect 193306 518058 193542 518294
rect 199826 705562 200062 705798
rect 200146 705562 200382 705798
rect 199826 705242 200062 705478
rect 200146 705242 200382 705478
rect 199826 669218 200062 669454
rect 200146 669218 200382 669454
rect 199826 668898 200062 669134
rect 200146 668898 200382 669134
rect 199826 633218 200062 633454
rect 200146 633218 200382 633454
rect 199826 632898 200062 633134
rect 200146 632898 200382 633134
rect 199826 597218 200062 597454
rect 200146 597218 200382 597454
rect 199826 596898 200062 597134
rect 200146 596898 200382 597134
rect 199826 561218 200062 561454
rect 200146 561218 200382 561454
rect 199826 560898 200062 561134
rect 200146 560898 200382 561134
rect 199826 525218 200062 525454
rect 200146 525218 200382 525454
rect 199826 524898 200062 525134
rect 200146 524898 200382 525134
rect 203546 672938 203782 673174
rect 203866 672938 204102 673174
rect 203546 672618 203782 672854
rect 203866 672618 204102 672854
rect 203546 636938 203782 637174
rect 203866 636938 204102 637174
rect 203546 636618 203782 636854
rect 203866 636618 204102 636854
rect 203546 600938 203782 601174
rect 203866 600938 204102 601174
rect 203546 600618 203782 600854
rect 203866 600618 204102 600854
rect 203546 564938 203782 565174
rect 203866 564938 204102 565174
rect 203546 564618 203782 564854
rect 203866 564618 204102 564854
rect 203546 528938 203782 529174
rect 203866 528938 204102 529174
rect 203546 528618 203782 528854
rect 203866 528618 204102 528854
rect 207266 676658 207502 676894
rect 207586 676658 207822 676894
rect 207266 676338 207502 676574
rect 207586 676338 207822 676574
rect 207266 640658 207502 640894
rect 207586 640658 207822 640894
rect 207266 640338 207502 640574
rect 207586 640338 207822 640574
rect 207266 604658 207502 604894
rect 207586 604658 207822 604894
rect 207266 604338 207502 604574
rect 207586 604338 207822 604574
rect 207266 568658 207502 568894
rect 207586 568658 207822 568894
rect 207266 568338 207502 568574
rect 207586 568338 207822 568574
rect 207266 532658 207502 532894
rect 207586 532658 207822 532894
rect 207266 532338 207502 532574
rect 207586 532338 207822 532574
rect 228986 710362 229222 710598
rect 229306 710362 229542 710598
rect 228986 710042 229222 710278
rect 229306 710042 229542 710278
rect 225266 708442 225502 708678
rect 225586 708442 225822 708678
rect 225266 708122 225502 708358
rect 225586 708122 225822 708358
rect 221546 706522 221782 706758
rect 221866 706522 222102 706758
rect 221546 706202 221782 706438
rect 221866 706202 222102 706438
rect 210986 680378 211222 680614
rect 211306 680378 211542 680614
rect 210986 680058 211222 680294
rect 211306 680058 211542 680294
rect 210986 644378 211222 644614
rect 211306 644378 211542 644614
rect 210986 644058 211222 644294
rect 211306 644058 211542 644294
rect 210986 608378 211222 608614
rect 211306 608378 211542 608614
rect 210986 608058 211222 608294
rect 211306 608058 211542 608294
rect 210986 572378 211222 572614
rect 211306 572378 211542 572614
rect 210986 572058 211222 572294
rect 211306 572058 211542 572294
rect 210986 536378 211222 536614
rect 211306 536378 211542 536614
rect 210986 536058 211222 536294
rect 211306 536058 211542 536294
rect 217826 704602 218062 704838
rect 218146 704602 218382 704838
rect 217826 704282 218062 704518
rect 218146 704282 218382 704518
rect 217826 687218 218062 687454
rect 218146 687218 218382 687454
rect 217826 686898 218062 687134
rect 218146 686898 218382 687134
rect 217826 651218 218062 651454
rect 218146 651218 218382 651454
rect 217826 650898 218062 651134
rect 218146 650898 218382 651134
rect 217826 615218 218062 615454
rect 218146 615218 218382 615454
rect 217826 614898 218062 615134
rect 218146 614898 218382 615134
rect 217826 579218 218062 579454
rect 218146 579218 218382 579454
rect 217826 578898 218062 579134
rect 218146 578898 218382 579134
rect 217826 543218 218062 543454
rect 218146 543218 218382 543454
rect 217826 542898 218062 543134
rect 218146 542898 218382 543134
rect 221546 690938 221782 691174
rect 221866 690938 222102 691174
rect 221546 690618 221782 690854
rect 221866 690618 222102 690854
rect 221546 654938 221782 655174
rect 221866 654938 222102 655174
rect 221546 654618 221782 654854
rect 221866 654618 222102 654854
rect 221546 618938 221782 619174
rect 221866 618938 222102 619174
rect 221546 618618 221782 618854
rect 221866 618618 222102 618854
rect 221546 582938 221782 583174
rect 221866 582938 222102 583174
rect 221546 582618 221782 582854
rect 221866 582618 222102 582854
rect 221546 546938 221782 547174
rect 221866 546938 222102 547174
rect 221546 546618 221782 546854
rect 221866 546618 222102 546854
rect 221546 510938 221782 511174
rect 221866 510938 222102 511174
rect 221546 510618 221782 510854
rect 221866 510618 222102 510854
rect 225266 694658 225502 694894
rect 225586 694658 225822 694894
rect 225266 694338 225502 694574
rect 225586 694338 225822 694574
rect 225266 658658 225502 658894
rect 225586 658658 225822 658894
rect 225266 658338 225502 658574
rect 225586 658338 225822 658574
rect 225266 622658 225502 622894
rect 225586 622658 225822 622894
rect 225266 622338 225502 622574
rect 225586 622338 225822 622574
rect 225266 586658 225502 586894
rect 225586 586658 225822 586894
rect 225266 586338 225502 586574
rect 225586 586338 225822 586574
rect 225266 550658 225502 550894
rect 225586 550658 225822 550894
rect 225266 550338 225502 550574
rect 225586 550338 225822 550574
rect 225266 514658 225502 514894
rect 225586 514658 225822 514894
rect 225266 514338 225502 514574
rect 225586 514338 225822 514574
rect 246986 711322 247222 711558
rect 247306 711322 247542 711558
rect 246986 711002 247222 711238
rect 247306 711002 247542 711238
rect 243266 709402 243502 709638
rect 243586 709402 243822 709638
rect 243266 709082 243502 709318
rect 243586 709082 243822 709318
rect 239546 707482 239782 707718
rect 239866 707482 240102 707718
rect 239546 707162 239782 707398
rect 239866 707162 240102 707398
rect 228986 698378 229222 698614
rect 229306 698378 229542 698614
rect 228986 698058 229222 698294
rect 229306 698058 229542 698294
rect 228986 662378 229222 662614
rect 229306 662378 229542 662614
rect 228986 662058 229222 662294
rect 229306 662058 229542 662294
rect 228986 626378 229222 626614
rect 229306 626378 229542 626614
rect 228986 626058 229222 626294
rect 229306 626058 229542 626294
rect 228986 590378 229222 590614
rect 229306 590378 229542 590614
rect 228986 590058 229222 590294
rect 229306 590058 229542 590294
rect 228986 554378 229222 554614
rect 229306 554378 229542 554614
rect 228986 554058 229222 554294
rect 229306 554058 229542 554294
rect 228986 518378 229222 518614
rect 229306 518378 229542 518614
rect 228986 518058 229222 518294
rect 229306 518058 229542 518294
rect 235826 705562 236062 705798
rect 236146 705562 236382 705798
rect 235826 705242 236062 705478
rect 236146 705242 236382 705478
rect 235826 669218 236062 669454
rect 236146 669218 236382 669454
rect 235826 668898 236062 669134
rect 236146 668898 236382 669134
rect 235826 633218 236062 633454
rect 236146 633218 236382 633454
rect 235826 632898 236062 633134
rect 236146 632898 236382 633134
rect 235826 597218 236062 597454
rect 236146 597218 236382 597454
rect 235826 596898 236062 597134
rect 236146 596898 236382 597134
rect 235826 561218 236062 561454
rect 236146 561218 236382 561454
rect 235826 560898 236062 561134
rect 236146 560898 236382 561134
rect 235826 525218 236062 525454
rect 236146 525218 236382 525454
rect 235826 524898 236062 525134
rect 236146 524898 236382 525134
rect 239546 672938 239782 673174
rect 239866 672938 240102 673174
rect 239546 672618 239782 672854
rect 239866 672618 240102 672854
rect 239546 636938 239782 637174
rect 239866 636938 240102 637174
rect 239546 636618 239782 636854
rect 239866 636618 240102 636854
rect 239546 600938 239782 601174
rect 239866 600938 240102 601174
rect 239546 600618 239782 600854
rect 239866 600618 240102 600854
rect 239546 564938 239782 565174
rect 239866 564938 240102 565174
rect 239546 564618 239782 564854
rect 239866 564618 240102 564854
rect 239546 528938 239782 529174
rect 239866 528938 240102 529174
rect 239546 528618 239782 528854
rect 239866 528618 240102 528854
rect 243266 676658 243502 676894
rect 243586 676658 243822 676894
rect 243266 676338 243502 676574
rect 243586 676338 243822 676574
rect 243266 640658 243502 640894
rect 243586 640658 243822 640894
rect 243266 640338 243502 640574
rect 243586 640338 243822 640574
rect 243266 604658 243502 604894
rect 243586 604658 243822 604894
rect 243266 604338 243502 604574
rect 243586 604338 243822 604574
rect 243266 568658 243502 568894
rect 243586 568658 243822 568894
rect 243266 568338 243502 568574
rect 243586 568338 243822 568574
rect 243266 532658 243502 532894
rect 243586 532658 243822 532894
rect 243266 532338 243502 532574
rect 243586 532338 243822 532574
rect 264986 710362 265222 710598
rect 265306 710362 265542 710598
rect 264986 710042 265222 710278
rect 265306 710042 265542 710278
rect 261266 708442 261502 708678
rect 261586 708442 261822 708678
rect 261266 708122 261502 708358
rect 261586 708122 261822 708358
rect 257546 706522 257782 706758
rect 257866 706522 258102 706758
rect 257546 706202 257782 706438
rect 257866 706202 258102 706438
rect 246986 680378 247222 680614
rect 247306 680378 247542 680614
rect 246986 680058 247222 680294
rect 247306 680058 247542 680294
rect 246986 644378 247222 644614
rect 247306 644378 247542 644614
rect 246986 644058 247222 644294
rect 247306 644058 247542 644294
rect 246986 608378 247222 608614
rect 247306 608378 247542 608614
rect 246986 608058 247222 608294
rect 247306 608058 247542 608294
rect 246986 572378 247222 572614
rect 247306 572378 247542 572614
rect 246986 572058 247222 572294
rect 247306 572058 247542 572294
rect 246986 536378 247222 536614
rect 247306 536378 247542 536614
rect 246986 536058 247222 536294
rect 247306 536058 247542 536294
rect 253826 704602 254062 704838
rect 254146 704602 254382 704838
rect 253826 704282 254062 704518
rect 254146 704282 254382 704518
rect 253826 687218 254062 687454
rect 254146 687218 254382 687454
rect 253826 686898 254062 687134
rect 254146 686898 254382 687134
rect 253826 651218 254062 651454
rect 254146 651218 254382 651454
rect 253826 650898 254062 651134
rect 254146 650898 254382 651134
rect 253826 615218 254062 615454
rect 254146 615218 254382 615454
rect 253826 614898 254062 615134
rect 254146 614898 254382 615134
rect 253826 579218 254062 579454
rect 254146 579218 254382 579454
rect 253826 578898 254062 579134
rect 254146 578898 254382 579134
rect 253826 543218 254062 543454
rect 254146 543218 254382 543454
rect 253826 542898 254062 543134
rect 254146 542898 254382 543134
rect 257546 690938 257782 691174
rect 257866 690938 258102 691174
rect 257546 690618 257782 690854
rect 257866 690618 258102 690854
rect 257546 654938 257782 655174
rect 257866 654938 258102 655174
rect 257546 654618 257782 654854
rect 257866 654618 258102 654854
rect 257546 618938 257782 619174
rect 257866 618938 258102 619174
rect 257546 618618 257782 618854
rect 257866 618618 258102 618854
rect 257546 582938 257782 583174
rect 257866 582938 258102 583174
rect 257546 582618 257782 582854
rect 257866 582618 258102 582854
rect 257546 546938 257782 547174
rect 257866 546938 258102 547174
rect 257546 546618 257782 546854
rect 257866 546618 258102 546854
rect 257546 510938 257782 511174
rect 257866 510938 258102 511174
rect 257546 510618 257782 510854
rect 257866 510618 258102 510854
rect 261266 694658 261502 694894
rect 261586 694658 261822 694894
rect 261266 694338 261502 694574
rect 261586 694338 261822 694574
rect 261266 658658 261502 658894
rect 261586 658658 261822 658894
rect 261266 658338 261502 658574
rect 261586 658338 261822 658574
rect 261266 622658 261502 622894
rect 261586 622658 261822 622894
rect 261266 622338 261502 622574
rect 261586 622338 261822 622574
rect 261266 586658 261502 586894
rect 261586 586658 261822 586894
rect 261266 586338 261502 586574
rect 261586 586338 261822 586574
rect 261266 550658 261502 550894
rect 261586 550658 261822 550894
rect 261266 550338 261502 550574
rect 261586 550338 261822 550574
rect 261266 514658 261502 514894
rect 261586 514658 261822 514894
rect 261266 514338 261502 514574
rect 261586 514338 261822 514574
rect 282986 711322 283222 711558
rect 283306 711322 283542 711558
rect 282986 711002 283222 711238
rect 283306 711002 283542 711238
rect 279266 709402 279502 709638
rect 279586 709402 279822 709638
rect 279266 709082 279502 709318
rect 279586 709082 279822 709318
rect 275546 707482 275782 707718
rect 275866 707482 276102 707718
rect 275546 707162 275782 707398
rect 275866 707162 276102 707398
rect 264986 698378 265222 698614
rect 265306 698378 265542 698614
rect 264986 698058 265222 698294
rect 265306 698058 265542 698294
rect 264986 662378 265222 662614
rect 265306 662378 265542 662614
rect 264986 662058 265222 662294
rect 265306 662058 265542 662294
rect 264986 626378 265222 626614
rect 265306 626378 265542 626614
rect 264986 626058 265222 626294
rect 265306 626058 265542 626294
rect 264986 590378 265222 590614
rect 265306 590378 265542 590614
rect 264986 590058 265222 590294
rect 265306 590058 265542 590294
rect 264986 554378 265222 554614
rect 265306 554378 265542 554614
rect 264986 554058 265222 554294
rect 265306 554058 265542 554294
rect 264986 518378 265222 518614
rect 265306 518378 265542 518614
rect 264986 518058 265222 518294
rect 265306 518058 265542 518294
rect 271826 705562 272062 705798
rect 272146 705562 272382 705798
rect 271826 705242 272062 705478
rect 272146 705242 272382 705478
rect 271826 669218 272062 669454
rect 272146 669218 272382 669454
rect 271826 668898 272062 669134
rect 272146 668898 272382 669134
rect 271826 633218 272062 633454
rect 272146 633218 272382 633454
rect 271826 632898 272062 633134
rect 272146 632898 272382 633134
rect 271826 597218 272062 597454
rect 272146 597218 272382 597454
rect 271826 596898 272062 597134
rect 272146 596898 272382 597134
rect 271826 561218 272062 561454
rect 272146 561218 272382 561454
rect 271826 560898 272062 561134
rect 272146 560898 272382 561134
rect 271826 525218 272062 525454
rect 272146 525218 272382 525454
rect 271826 524898 272062 525134
rect 272146 524898 272382 525134
rect 275546 672938 275782 673174
rect 275866 672938 276102 673174
rect 275546 672618 275782 672854
rect 275866 672618 276102 672854
rect 275546 636938 275782 637174
rect 275866 636938 276102 637174
rect 275546 636618 275782 636854
rect 275866 636618 276102 636854
rect 275546 600938 275782 601174
rect 275866 600938 276102 601174
rect 275546 600618 275782 600854
rect 275866 600618 276102 600854
rect 275546 564938 275782 565174
rect 275866 564938 276102 565174
rect 275546 564618 275782 564854
rect 275866 564618 276102 564854
rect 275546 528938 275782 529174
rect 275866 528938 276102 529174
rect 275546 528618 275782 528854
rect 275866 528618 276102 528854
rect 279266 676658 279502 676894
rect 279586 676658 279822 676894
rect 279266 676338 279502 676574
rect 279586 676338 279822 676574
rect 279266 640658 279502 640894
rect 279586 640658 279822 640894
rect 279266 640338 279502 640574
rect 279586 640338 279822 640574
rect 279266 604658 279502 604894
rect 279586 604658 279822 604894
rect 279266 604338 279502 604574
rect 279586 604338 279822 604574
rect 279266 568658 279502 568894
rect 279586 568658 279822 568894
rect 279266 568338 279502 568574
rect 279586 568338 279822 568574
rect 279266 532658 279502 532894
rect 279586 532658 279822 532894
rect 279266 532338 279502 532574
rect 279586 532338 279822 532574
rect 300986 710362 301222 710598
rect 301306 710362 301542 710598
rect 300986 710042 301222 710278
rect 301306 710042 301542 710278
rect 297266 708442 297502 708678
rect 297586 708442 297822 708678
rect 297266 708122 297502 708358
rect 297586 708122 297822 708358
rect 293546 706522 293782 706758
rect 293866 706522 294102 706758
rect 293546 706202 293782 706438
rect 293866 706202 294102 706438
rect 282986 680378 283222 680614
rect 283306 680378 283542 680614
rect 282986 680058 283222 680294
rect 283306 680058 283542 680294
rect 282986 644378 283222 644614
rect 283306 644378 283542 644614
rect 282986 644058 283222 644294
rect 283306 644058 283542 644294
rect 282986 608378 283222 608614
rect 283306 608378 283542 608614
rect 282986 608058 283222 608294
rect 283306 608058 283542 608294
rect 282986 572378 283222 572614
rect 283306 572378 283542 572614
rect 282986 572058 283222 572294
rect 283306 572058 283542 572294
rect 282986 536378 283222 536614
rect 283306 536378 283542 536614
rect 282986 536058 283222 536294
rect 283306 536058 283542 536294
rect 289826 704602 290062 704838
rect 290146 704602 290382 704838
rect 289826 704282 290062 704518
rect 290146 704282 290382 704518
rect 289826 687218 290062 687454
rect 290146 687218 290382 687454
rect 289826 686898 290062 687134
rect 290146 686898 290382 687134
rect 289826 651218 290062 651454
rect 290146 651218 290382 651454
rect 289826 650898 290062 651134
rect 290146 650898 290382 651134
rect 289826 615218 290062 615454
rect 290146 615218 290382 615454
rect 289826 614898 290062 615134
rect 290146 614898 290382 615134
rect 289826 579218 290062 579454
rect 290146 579218 290382 579454
rect 289826 578898 290062 579134
rect 290146 578898 290382 579134
rect 289826 543218 290062 543454
rect 290146 543218 290382 543454
rect 289826 542898 290062 543134
rect 290146 542898 290382 543134
rect 293546 690938 293782 691174
rect 293866 690938 294102 691174
rect 293546 690618 293782 690854
rect 293866 690618 294102 690854
rect 293546 654938 293782 655174
rect 293866 654938 294102 655174
rect 293546 654618 293782 654854
rect 293866 654618 294102 654854
rect 293546 618938 293782 619174
rect 293866 618938 294102 619174
rect 293546 618618 293782 618854
rect 293866 618618 294102 618854
rect 293546 582938 293782 583174
rect 293866 582938 294102 583174
rect 293546 582618 293782 582854
rect 293866 582618 294102 582854
rect 293546 546938 293782 547174
rect 293866 546938 294102 547174
rect 293546 546618 293782 546854
rect 293866 546618 294102 546854
rect 293546 510938 293782 511174
rect 293866 510938 294102 511174
rect 293546 510618 293782 510854
rect 293866 510618 294102 510854
rect 297266 694658 297502 694894
rect 297586 694658 297822 694894
rect 297266 694338 297502 694574
rect 297586 694338 297822 694574
rect 297266 658658 297502 658894
rect 297586 658658 297822 658894
rect 297266 658338 297502 658574
rect 297586 658338 297822 658574
rect 297266 622658 297502 622894
rect 297586 622658 297822 622894
rect 297266 622338 297502 622574
rect 297586 622338 297822 622574
rect 297266 586658 297502 586894
rect 297586 586658 297822 586894
rect 297266 586338 297502 586574
rect 297586 586338 297822 586574
rect 297266 550658 297502 550894
rect 297586 550658 297822 550894
rect 297266 550338 297502 550574
rect 297586 550338 297822 550574
rect 297266 514658 297502 514894
rect 297586 514658 297822 514894
rect 297266 514338 297502 514574
rect 297586 514338 297822 514574
rect 318986 711322 319222 711558
rect 319306 711322 319542 711558
rect 318986 711002 319222 711238
rect 319306 711002 319542 711238
rect 315266 709402 315502 709638
rect 315586 709402 315822 709638
rect 315266 709082 315502 709318
rect 315586 709082 315822 709318
rect 311546 707482 311782 707718
rect 311866 707482 312102 707718
rect 311546 707162 311782 707398
rect 311866 707162 312102 707398
rect 300986 698378 301222 698614
rect 301306 698378 301542 698614
rect 300986 698058 301222 698294
rect 301306 698058 301542 698294
rect 300986 662378 301222 662614
rect 301306 662378 301542 662614
rect 300986 662058 301222 662294
rect 301306 662058 301542 662294
rect 300986 626378 301222 626614
rect 301306 626378 301542 626614
rect 300986 626058 301222 626294
rect 301306 626058 301542 626294
rect 300986 590378 301222 590614
rect 301306 590378 301542 590614
rect 300986 590058 301222 590294
rect 301306 590058 301542 590294
rect 300986 554378 301222 554614
rect 301306 554378 301542 554614
rect 300986 554058 301222 554294
rect 301306 554058 301542 554294
rect 300986 518378 301222 518614
rect 301306 518378 301542 518614
rect 300986 518058 301222 518294
rect 301306 518058 301542 518294
rect 307826 705562 308062 705798
rect 308146 705562 308382 705798
rect 307826 705242 308062 705478
rect 308146 705242 308382 705478
rect 307826 669218 308062 669454
rect 308146 669218 308382 669454
rect 307826 668898 308062 669134
rect 308146 668898 308382 669134
rect 307826 633218 308062 633454
rect 308146 633218 308382 633454
rect 307826 632898 308062 633134
rect 308146 632898 308382 633134
rect 307826 597218 308062 597454
rect 308146 597218 308382 597454
rect 307826 596898 308062 597134
rect 308146 596898 308382 597134
rect 307826 561218 308062 561454
rect 308146 561218 308382 561454
rect 307826 560898 308062 561134
rect 308146 560898 308382 561134
rect 307826 525218 308062 525454
rect 308146 525218 308382 525454
rect 307826 524898 308062 525134
rect 308146 524898 308382 525134
rect 311546 672938 311782 673174
rect 311866 672938 312102 673174
rect 311546 672618 311782 672854
rect 311866 672618 312102 672854
rect 311546 636938 311782 637174
rect 311866 636938 312102 637174
rect 311546 636618 311782 636854
rect 311866 636618 312102 636854
rect 311546 600938 311782 601174
rect 311866 600938 312102 601174
rect 311546 600618 311782 600854
rect 311866 600618 312102 600854
rect 311546 564938 311782 565174
rect 311866 564938 312102 565174
rect 311546 564618 311782 564854
rect 311866 564618 312102 564854
rect 311546 528938 311782 529174
rect 311866 528938 312102 529174
rect 311546 528618 311782 528854
rect 311866 528618 312102 528854
rect 315266 676658 315502 676894
rect 315586 676658 315822 676894
rect 315266 676338 315502 676574
rect 315586 676338 315822 676574
rect 315266 640658 315502 640894
rect 315586 640658 315822 640894
rect 315266 640338 315502 640574
rect 315586 640338 315822 640574
rect 315266 604658 315502 604894
rect 315586 604658 315822 604894
rect 315266 604338 315502 604574
rect 315586 604338 315822 604574
rect 315266 568658 315502 568894
rect 315586 568658 315822 568894
rect 315266 568338 315502 568574
rect 315586 568338 315822 568574
rect 315266 532658 315502 532894
rect 315586 532658 315822 532894
rect 315266 532338 315502 532574
rect 315586 532338 315822 532574
rect 336986 710362 337222 710598
rect 337306 710362 337542 710598
rect 336986 710042 337222 710278
rect 337306 710042 337542 710278
rect 333266 708442 333502 708678
rect 333586 708442 333822 708678
rect 333266 708122 333502 708358
rect 333586 708122 333822 708358
rect 329546 706522 329782 706758
rect 329866 706522 330102 706758
rect 329546 706202 329782 706438
rect 329866 706202 330102 706438
rect 318986 680378 319222 680614
rect 319306 680378 319542 680614
rect 318986 680058 319222 680294
rect 319306 680058 319542 680294
rect 318986 644378 319222 644614
rect 319306 644378 319542 644614
rect 318986 644058 319222 644294
rect 319306 644058 319542 644294
rect 318986 608378 319222 608614
rect 319306 608378 319542 608614
rect 318986 608058 319222 608294
rect 319306 608058 319542 608294
rect 318986 572378 319222 572614
rect 319306 572378 319542 572614
rect 318986 572058 319222 572294
rect 319306 572058 319542 572294
rect 318986 536378 319222 536614
rect 319306 536378 319542 536614
rect 318986 536058 319222 536294
rect 319306 536058 319542 536294
rect 325826 704602 326062 704838
rect 326146 704602 326382 704838
rect 325826 704282 326062 704518
rect 326146 704282 326382 704518
rect 325826 687218 326062 687454
rect 326146 687218 326382 687454
rect 325826 686898 326062 687134
rect 326146 686898 326382 687134
rect 325826 651218 326062 651454
rect 326146 651218 326382 651454
rect 325826 650898 326062 651134
rect 326146 650898 326382 651134
rect 325826 615218 326062 615454
rect 326146 615218 326382 615454
rect 325826 614898 326062 615134
rect 326146 614898 326382 615134
rect 325826 579218 326062 579454
rect 326146 579218 326382 579454
rect 325826 578898 326062 579134
rect 326146 578898 326382 579134
rect 325826 543218 326062 543454
rect 326146 543218 326382 543454
rect 325826 542898 326062 543134
rect 326146 542898 326382 543134
rect 329546 690938 329782 691174
rect 329866 690938 330102 691174
rect 329546 690618 329782 690854
rect 329866 690618 330102 690854
rect 329546 654938 329782 655174
rect 329866 654938 330102 655174
rect 329546 654618 329782 654854
rect 329866 654618 330102 654854
rect 329546 618938 329782 619174
rect 329866 618938 330102 619174
rect 329546 618618 329782 618854
rect 329866 618618 330102 618854
rect 329546 582938 329782 583174
rect 329866 582938 330102 583174
rect 329546 582618 329782 582854
rect 329866 582618 330102 582854
rect 329546 546938 329782 547174
rect 329866 546938 330102 547174
rect 329546 546618 329782 546854
rect 329866 546618 330102 546854
rect 329546 510938 329782 511174
rect 329866 510938 330102 511174
rect 329546 510618 329782 510854
rect 329866 510618 330102 510854
rect 333266 694658 333502 694894
rect 333586 694658 333822 694894
rect 333266 694338 333502 694574
rect 333586 694338 333822 694574
rect 333266 658658 333502 658894
rect 333586 658658 333822 658894
rect 333266 658338 333502 658574
rect 333586 658338 333822 658574
rect 333266 622658 333502 622894
rect 333586 622658 333822 622894
rect 333266 622338 333502 622574
rect 333586 622338 333822 622574
rect 333266 586658 333502 586894
rect 333586 586658 333822 586894
rect 333266 586338 333502 586574
rect 333586 586338 333822 586574
rect 333266 550658 333502 550894
rect 333586 550658 333822 550894
rect 333266 550338 333502 550574
rect 333586 550338 333822 550574
rect 333266 514658 333502 514894
rect 333586 514658 333822 514894
rect 333266 514338 333502 514574
rect 333586 514338 333822 514574
rect 354986 711322 355222 711558
rect 355306 711322 355542 711558
rect 354986 711002 355222 711238
rect 355306 711002 355542 711238
rect 351266 709402 351502 709638
rect 351586 709402 351822 709638
rect 351266 709082 351502 709318
rect 351586 709082 351822 709318
rect 347546 707482 347782 707718
rect 347866 707482 348102 707718
rect 347546 707162 347782 707398
rect 347866 707162 348102 707398
rect 336986 698378 337222 698614
rect 337306 698378 337542 698614
rect 336986 698058 337222 698294
rect 337306 698058 337542 698294
rect 336986 662378 337222 662614
rect 337306 662378 337542 662614
rect 336986 662058 337222 662294
rect 337306 662058 337542 662294
rect 336986 626378 337222 626614
rect 337306 626378 337542 626614
rect 336986 626058 337222 626294
rect 337306 626058 337542 626294
rect 336986 590378 337222 590614
rect 337306 590378 337542 590614
rect 336986 590058 337222 590294
rect 337306 590058 337542 590294
rect 336986 554378 337222 554614
rect 337306 554378 337542 554614
rect 336986 554058 337222 554294
rect 337306 554058 337542 554294
rect 336986 518378 337222 518614
rect 337306 518378 337542 518614
rect 336986 518058 337222 518294
rect 337306 518058 337542 518294
rect 343826 705562 344062 705798
rect 344146 705562 344382 705798
rect 343826 705242 344062 705478
rect 344146 705242 344382 705478
rect 343826 669218 344062 669454
rect 344146 669218 344382 669454
rect 343826 668898 344062 669134
rect 344146 668898 344382 669134
rect 343826 633218 344062 633454
rect 344146 633218 344382 633454
rect 343826 632898 344062 633134
rect 344146 632898 344382 633134
rect 343826 597218 344062 597454
rect 344146 597218 344382 597454
rect 343826 596898 344062 597134
rect 344146 596898 344382 597134
rect 343826 561218 344062 561454
rect 344146 561218 344382 561454
rect 343826 560898 344062 561134
rect 344146 560898 344382 561134
rect 343826 525218 344062 525454
rect 344146 525218 344382 525454
rect 343826 524898 344062 525134
rect 344146 524898 344382 525134
rect 347546 672938 347782 673174
rect 347866 672938 348102 673174
rect 347546 672618 347782 672854
rect 347866 672618 348102 672854
rect 347546 636938 347782 637174
rect 347866 636938 348102 637174
rect 347546 636618 347782 636854
rect 347866 636618 348102 636854
rect 347546 600938 347782 601174
rect 347866 600938 348102 601174
rect 347546 600618 347782 600854
rect 347866 600618 348102 600854
rect 347546 564938 347782 565174
rect 347866 564938 348102 565174
rect 347546 564618 347782 564854
rect 347866 564618 348102 564854
rect 347546 528938 347782 529174
rect 347866 528938 348102 529174
rect 347546 528618 347782 528854
rect 347866 528618 348102 528854
rect 351266 676658 351502 676894
rect 351586 676658 351822 676894
rect 351266 676338 351502 676574
rect 351586 676338 351822 676574
rect 351266 640658 351502 640894
rect 351586 640658 351822 640894
rect 351266 640338 351502 640574
rect 351586 640338 351822 640574
rect 351266 604658 351502 604894
rect 351586 604658 351822 604894
rect 351266 604338 351502 604574
rect 351586 604338 351822 604574
rect 351266 568658 351502 568894
rect 351586 568658 351822 568894
rect 351266 568338 351502 568574
rect 351586 568338 351822 568574
rect 351266 532658 351502 532894
rect 351586 532658 351822 532894
rect 351266 532338 351502 532574
rect 351586 532338 351822 532574
rect 372986 710362 373222 710598
rect 373306 710362 373542 710598
rect 372986 710042 373222 710278
rect 373306 710042 373542 710278
rect 369266 708442 369502 708678
rect 369586 708442 369822 708678
rect 369266 708122 369502 708358
rect 369586 708122 369822 708358
rect 365546 706522 365782 706758
rect 365866 706522 366102 706758
rect 365546 706202 365782 706438
rect 365866 706202 366102 706438
rect 354986 680378 355222 680614
rect 355306 680378 355542 680614
rect 354986 680058 355222 680294
rect 355306 680058 355542 680294
rect 354986 644378 355222 644614
rect 355306 644378 355542 644614
rect 354986 644058 355222 644294
rect 355306 644058 355542 644294
rect 354986 608378 355222 608614
rect 355306 608378 355542 608614
rect 354986 608058 355222 608294
rect 355306 608058 355542 608294
rect 354986 572378 355222 572614
rect 355306 572378 355542 572614
rect 354986 572058 355222 572294
rect 355306 572058 355542 572294
rect 354986 536378 355222 536614
rect 355306 536378 355542 536614
rect 354986 536058 355222 536294
rect 355306 536058 355542 536294
rect 361826 704602 362062 704838
rect 362146 704602 362382 704838
rect 361826 704282 362062 704518
rect 362146 704282 362382 704518
rect 361826 687218 362062 687454
rect 362146 687218 362382 687454
rect 361826 686898 362062 687134
rect 362146 686898 362382 687134
rect 361826 651218 362062 651454
rect 362146 651218 362382 651454
rect 361826 650898 362062 651134
rect 362146 650898 362382 651134
rect 361826 615218 362062 615454
rect 362146 615218 362382 615454
rect 361826 614898 362062 615134
rect 362146 614898 362382 615134
rect 361826 579218 362062 579454
rect 362146 579218 362382 579454
rect 361826 578898 362062 579134
rect 362146 578898 362382 579134
rect 361826 543218 362062 543454
rect 362146 543218 362382 543454
rect 361826 542898 362062 543134
rect 362146 542898 362382 543134
rect 365546 690938 365782 691174
rect 365866 690938 366102 691174
rect 365546 690618 365782 690854
rect 365866 690618 366102 690854
rect 365546 654938 365782 655174
rect 365866 654938 366102 655174
rect 365546 654618 365782 654854
rect 365866 654618 366102 654854
rect 365546 618938 365782 619174
rect 365866 618938 366102 619174
rect 365546 618618 365782 618854
rect 365866 618618 366102 618854
rect 365546 582938 365782 583174
rect 365866 582938 366102 583174
rect 365546 582618 365782 582854
rect 365866 582618 366102 582854
rect 365546 546938 365782 547174
rect 365866 546938 366102 547174
rect 365546 546618 365782 546854
rect 365866 546618 366102 546854
rect 365546 510938 365782 511174
rect 365866 510938 366102 511174
rect 365546 510618 365782 510854
rect 365866 510618 366102 510854
rect 369266 694658 369502 694894
rect 369586 694658 369822 694894
rect 369266 694338 369502 694574
rect 369586 694338 369822 694574
rect 369266 658658 369502 658894
rect 369586 658658 369822 658894
rect 369266 658338 369502 658574
rect 369586 658338 369822 658574
rect 369266 622658 369502 622894
rect 369586 622658 369822 622894
rect 369266 622338 369502 622574
rect 369586 622338 369822 622574
rect 369266 586658 369502 586894
rect 369586 586658 369822 586894
rect 369266 586338 369502 586574
rect 369586 586338 369822 586574
rect 369266 550658 369502 550894
rect 369586 550658 369822 550894
rect 369266 550338 369502 550574
rect 369586 550338 369822 550574
rect 369266 514658 369502 514894
rect 369586 514658 369822 514894
rect 369266 514338 369502 514574
rect 369586 514338 369822 514574
rect 390986 711322 391222 711558
rect 391306 711322 391542 711558
rect 390986 711002 391222 711238
rect 391306 711002 391542 711238
rect 387266 709402 387502 709638
rect 387586 709402 387822 709638
rect 387266 709082 387502 709318
rect 387586 709082 387822 709318
rect 383546 707482 383782 707718
rect 383866 707482 384102 707718
rect 383546 707162 383782 707398
rect 383866 707162 384102 707398
rect 372986 698378 373222 698614
rect 373306 698378 373542 698614
rect 372986 698058 373222 698294
rect 373306 698058 373542 698294
rect 372986 662378 373222 662614
rect 373306 662378 373542 662614
rect 372986 662058 373222 662294
rect 373306 662058 373542 662294
rect 372986 626378 373222 626614
rect 373306 626378 373542 626614
rect 372986 626058 373222 626294
rect 373306 626058 373542 626294
rect 372986 590378 373222 590614
rect 373306 590378 373542 590614
rect 372986 590058 373222 590294
rect 373306 590058 373542 590294
rect 372986 554378 373222 554614
rect 373306 554378 373542 554614
rect 372986 554058 373222 554294
rect 373306 554058 373542 554294
rect 372986 518378 373222 518614
rect 373306 518378 373542 518614
rect 372986 518058 373222 518294
rect 373306 518058 373542 518294
rect 379826 705562 380062 705798
rect 380146 705562 380382 705798
rect 379826 705242 380062 705478
rect 380146 705242 380382 705478
rect 379826 669218 380062 669454
rect 380146 669218 380382 669454
rect 379826 668898 380062 669134
rect 380146 668898 380382 669134
rect 379826 633218 380062 633454
rect 380146 633218 380382 633454
rect 379826 632898 380062 633134
rect 380146 632898 380382 633134
rect 379826 597218 380062 597454
rect 380146 597218 380382 597454
rect 379826 596898 380062 597134
rect 380146 596898 380382 597134
rect 379826 561218 380062 561454
rect 380146 561218 380382 561454
rect 379826 560898 380062 561134
rect 380146 560898 380382 561134
rect 379826 525218 380062 525454
rect 380146 525218 380382 525454
rect 379826 524898 380062 525134
rect 380146 524898 380382 525134
rect 383546 672938 383782 673174
rect 383866 672938 384102 673174
rect 383546 672618 383782 672854
rect 383866 672618 384102 672854
rect 383546 636938 383782 637174
rect 383866 636938 384102 637174
rect 383546 636618 383782 636854
rect 383866 636618 384102 636854
rect 383546 600938 383782 601174
rect 383866 600938 384102 601174
rect 383546 600618 383782 600854
rect 383866 600618 384102 600854
rect 383546 564938 383782 565174
rect 383866 564938 384102 565174
rect 383546 564618 383782 564854
rect 383866 564618 384102 564854
rect 383546 528938 383782 529174
rect 383866 528938 384102 529174
rect 383546 528618 383782 528854
rect 383866 528618 384102 528854
rect 387266 676658 387502 676894
rect 387586 676658 387822 676894
rect 387266 676338 387502 676574
rect 387586 676338 387822 676574
rect 387266 640658 387502 640894
rect 387586 640658 387822 640894
rect 387266 640338 387502 640574
rect 387586 640338 387822 640574
rect 387266 604658 387502 604894
rect 387586 604658 387822 604894
rect 387266 604338 387502 604574
rect 387586 604338 387822 604574
rect 387266 568658 387502 568894
rect 387586 568658 387822 568894
rect 387266 568338 387502 568574
rect 387586 568338 387822 568574
rect 387266 532658 387502 532894
rect 387586 532658 387822 532894
rect 387266 532338 387502 532574
rect 387586 532338 387822 532574
rect 408986 710362 409222 710598
rect 409306 710362 409542 710598
rect 408986 710042 409222 710278
rect 409306 710042 409542 710278
rect 405266 708442 405502 708678
rect 405586 708442 405822 708678
rect 405266 708122 405502 708358
rect 405586 708122 405822 708358
rect 401546 706522 401782 706758
rect 401866 706522 402102 706758
rect 401546 706202 401782 706438
rect 401866 706202 402102 706438
rect 390986 680378 391222 680614
rect 391306 680378 391542 680614
rect 390986 680058 391222 680294
rect 391306 680058 391542 680294
rect 390986 644378 391222 644614
rect 391306 644378 391542 644614
rect 390986 644058 391222 644294
rect 391306 644058 391542 644294
rect 390986 608378 391222 608614
rect 391306 608378 391542 608614
rect 390986 608058 391222 608294
rect 391306 608058 391542 608294
rect 390986 572378 391222 572614
rect 391306 572378 391542 572614
rect 390986 572058 391222 572294
rect 391306 572058 391542 572294
rect 390986 536378 391222 536614
rect 391306 536378 391542 536614
rect 390986 536058 391222 536294
rect 391306 536058 391542 536294
rect 397826 704602 398062 704838
rect 398146 704602 398382 704838
rect 397826 704282 398062 704518
rect 398146 704282 398382 704518
rect 397826 687218 398062 687454
rect 398146 687218 398382 687454
rect 397826 686898 398062 687134
rect 398146 686898 398382 687134
rect 397826 651218 398062 651454
rect 398146 651218 398382 651454
rect 397826 650898 398062 651134
rect 398146 650898 398382 651134
rect 397826 615218 398062 615454
rect 398146 615218 398382 615454
rect 397826 614898 398062 615134
rect 398146 614898 398382 615134
rect 397826 579218 398062 579454
rect 398146 579218 398382 579454
rect 397826 578898 398062 579134
rect 398146 578898 398382 579134
rect 397826 543218 398062 543454
rect 398146 543218 398382 543454
rect 397826 542898 398062 543134
rect 398146 542898 398382 543134
rect 401546 690938 401782 691174
rect 401866 690938 402102 691174
rect 401546 690618 401782 690854
rect 401866 690618 402102 690854
rect 401546 654938 401782 655174
rect 401866 654938 402102 655174
rect 401546 654618 401782 654854
rect 401866 654618 402102 654854
rect 401546 618938 401782 619174
rect 401866 618938 402102 619174
rect 401546 618618 401782 618854
rect 401866 618618 402102 618854
rect 401546 582938 401782 583174
rect 401866 582938 402102 583174
rect 401546 582618 401782 582854
rect 401866 582618 402102 582854
rect 401546 546938 401782 547174
rect 401866 546938 402102 547174
rect 401546 546618 401782 546854
rect 401866 546618 402102 546854
rect 401546 510938 401782 511174
rect 401866 510938 402102 511174
rect 401546 510618 401782 510854
rect 401866 510618 402102 510854
rect 405266 694658 405502 694894
rect 405586 694658 405822 694894
rect 405266 694338 405502 694574
rect 405586 694338 405822 694574
rect 405266 658658 405502 658894
rect 405586 658658 405822 658894
rect 405266 658338 405502 658574
rect 405586 658338 405822 658574
rect 405266 622658 405502 622894
rect 405586 622658 405822 622894
rect 405266 622338 405502 622574
rect 405586 622338 405822 622574
rect 405266 586658 405502 586894
rect 405586 586658 405822 586894
rect 405266 586338 405502 586574
rect 405586 586338 405822 586574
rect 405266 550658 405502 550894
rect 405586 550658 405822 550894
rect 405266 550338 405502 550574
rect 405586 550338 405822 550574
rect 405266 514658 405502 514894
rect 405586 514658 405822 514894
rect 405266 514338 405502 514574
rect 405586 514338 405822 514574
rect 426986 711322 427222 711558
rect 427306 711322 427542 711558
rect 426986 711002 427222 711238
rect 427306 711002 427542 711238
rect 423266 709402 423502 709638
rect 423586 709402 423822 709638
rect 423266 709082 423502 709318
rect 423586 709082 423822 709318
rect 419546 707482 419782 707718
rect 419866 707482 420102 707718
rect 419546 707162 419782 707398
rect 419866 707162 420102 707398
rect 408986 698378 409222 698614
rect 409306 698378 409542 698614
rect 408986 698058 409222 698294
rect 409306 698058 409542 698294
rect 408986 662378 409222 662614
rect 409306 662378 409542 662614
rect 408986 662058 409222 662294
rect 409306 662058 409542 662294
rect 408986 626378 409222 626614
rect 409306 626378 409542 626614
rect 408986 626058 409222 626294
rect 409306 626058 409542 626294
rect 408986 590378 409222 590614
rect 409306 590378 409542 590614
rect 408986 590058 409222 590294
rect 409306 590058 409542 590294
rect 408986 554378 409222 554614
rect 409306 554378 409542 554614
rect 408986 554058 409222 554294
rect 409306 554058 409542 554294
rect 408986 518378 409222 518614
rect 409306 518378 409542 518614
rect 408986 518058 409222 518294
rect 409306 518058 409542 518294
rect 415826 705562 416062 705798
rect 416146 705562 416382 705798
rect 415826 705242 416062 705478
rect 416146 705242 416382 705478
rect 415826 669218 416062 669454
rect 416146 669218 416382 669454
rect 415826 668898 416062 669134
rect 416146 668898 416382 669134
rect 415826 633218 416062 633454
rect 416146 633218 416382 633454
rect 415826 632898 416062 633134
rect 416146 632898 416382 633134
rect 415826 597218 416062 597454
rect 416146 597218 416382 597454
rect 415826 596898 416062 597134
rect 416146 596898 416382 597134
rect 415826 561218 416062 561454
rect 416146 561218 416382 561454
rect 415826 560898 416062 561134
rect 416146 560898 416382 561134
rect 415826 525218 416062 525454
rect 416146 525218 416382 525454
rect 415826 524898 416062 525134
rect 416146 524898 416382 525134
rect 419546 672938 419782 673174
rect 419866 672938 420102 673174
rect 419546 672618 419782 672854
rect 419866 672618 420102 672854
rect 419546 636938 419782 637174
rect 419866 636938 420102 637174
rect 419546 636618 419782 636854
rect 419866 636618 420102 636854
rect 419546 600938 419782 601174
rect 419866 600938 420102 601174
rect 419546 600618 419782 600854
rect 419866 600618 420102 600854
rect 419546 564938 419782 565174
rect 419866 564938 420102 565174
rect 419546 564618 419782 564854
rect 419866 564618 420102 564854
rect 419546 528938 419782 529174
rect 419866 528938 420102 529174
rect 419546 528618 419782 528854
rect 419866 528618 420102 528854
rect 423266 676658 423502 676894
rect 423586 676658 423822 676894
rect 423266 676338 423502 676574
rect 423586 676338 423822 676574
rect 423266 640658 423502 640894
rect 423586 640658 423822 640894
rect 423266 640338 423502 640574
rect 423586 640338 423822 640574
rect 423266 604658 423502 604894
rect 423586 604658 423822 604894
rect 423266 604338 423502 604574
rect 423586 604338 423822 604574
rect 423266 568658 423502 568894
rect 423586 568658 423822 568894
rect 423266 568338 423502 568574
rect 423586 568338 423822 568574
rect 423266 532658 423502 532894
rect 423586 532658 423822 532894
rect 423266 532338 423502 532574
rect 423586 532338 423822 532574
rect 423266 496658 423502 496894
rect 423586 496658 423822 496894
rect 423266 496338 423502 496574
rect 423586 496338 423822 496574
rect 185410 489218 185646 489454
rect 185410 488898 185646 489134
rect 216130 489218 216366 489454
rect 216130 488898 216366 489134
rect 246850 489218 247086 489454
rect 246850 488898 247086 489134
rect 277570 489218 277806 489454
rect 277570 488898 277806 489134
rect 308290 489218 308526 489454
rect 308290 488898 308526 489134
rect 339010 489218 339246 489454
rect 339010 488898 339246 489134
rect 369730 489218 369966 489454
rect 369730 488898 369966 489134
rect 400450 489218 400686 489454
rect 400450 488898 400686 489134
rect 156986 482378 157222 482614
rect 157306 482378 157542 482614
rect 156986 482058 157222 482294
rect 157306 482058 157542 482294
rect 170050 471218 170286 471454
rect 170050 470898 170286 471134
rect 200770 471218 201006 471454
rect 200770 470898 201006 471134
rect 231490 471218 231726 471454
rect 231490 470898 231726 471134
rect 262210 471218 262446 471454
rect 262210 470898 262446 471134
rect 292930 471218 293166 471454
rect 292930 470898 293166 471134
rect 323650 471218 323886 471454
rect 323650 470898 323886 471134
rect 354370 471218 354606 471454
rect 354370 470898 354606 471134
rect 385090 471218 385326 471454
rect 385090 470898 385326 471134
rect 415810 471218 416046 471454
rect 415810 470898 416046 471134
rect 423266 460658 423502 460894
rect 423586 460658 423822 460894
rect 423266 460338 423502 460574
rect 423586 460338 423822 460574
rect 185410 453218 185646 453454
rect 185410 452898 185646 453134
rect 216130 453218 216366 453454
rect 216130 452898 216366 453134
rect 246850 453218 247086 453454
rect 246850 452898 247086 453134
rect 277570 453218 277806 453454
rect 277570 452898 277806 453134
rect 308290 453218 308526 453454
rect 308290 452898 308526 453134
rect 339010 453218 339246 453454
rect 339010 452898 339246 453134
rect 369730 453218 369966 453454
rect 369730 452898 369966 453134
rect 400450 453218 400686 453454
rect 400450 452898 400686 453134
rect 156986 446378 157222 446614
rect 157306 446378 157542 446614
rect 156986 446058 157222 446294
rect 157306 446058 157542 446294
rect 170050 435218 170286 435454
rect 170050 434898 170286 435134
rect 200770 435218 201006 435454
rect 200770 434898 201006 435134
rect 231490 435218 231726 435454
rect 231490 434898 231726 435134
rect 262210 435218 262446 435454
rect 262210 434898 262446 435134
rect 292930 435218 293166 435454
rect 292930 434898 293166 435134
rect 323650 435218 323886 435454
rect 323650 434898 323886 435134
rect 354370 435218 354606 435454
rect 354370 434898 354606 435134
rect 385090 435218 385326 435454
rect 385090 434898 385326 435134
rect 415810 435218 416046 435454
rect 415810 434898 416046 435134
rect 423266 424658 423502 424894
rect 423586 424658 423822 424894
rect 423266 424338 423502 424574
rect 423586 424338 423822 424574
rect 185410 417218 185646 417454
rect 185410 416898 185646 417134
rect 216130 417218 216366 417454
rect 216130 416898 216366 417134
rect 246850 417218 247086 417454
rect 246850 416898 247086 417134
rect 277570 417218 277806 417454
rect 277570 416898 277806 417134
rect 308290 417218 308526 417454
rect 308290 416898 308526 417134
rect 339010 417218 339246 417454
rect 339010 416898 339246 417134
rect 369730 417218 369966 417454
rect 369730 416898 369966 417134
rect 400450 417218 400686 417454
rect 400450 416898 400686 417134
rect 156986 410378 157222 410614
rect 157306 410378 157542 410614
rect 156986 410058 157222 410294
rect 157306 410058 157542 410294
rect 170050 399218 170286 399454
rect 170050 398898 170286 399134
rect 200770 399218 201006 399454
rect 200770 398898 201006 399134
rect 231490 399218 231726 399454
rect 231490 398898 231726 399134
rect 262210 399218 262446 399454
rect 262210 398898 262446 399134
rect 292930 399218 293166 399454
rect 292930 398898 293166 399134
rect 323650 399218 323886 399454
rect 323650 398898 323886 399134
rect 354370 399218 354606 399454
rect 354370 398898 354606 399134
rect 385090 399218 385326 399454
rect 385090 398898 385326 399134
rect 415810 399218 416046 399454
rect 415810 398898 416046 399134
rect 423266 388658 423502 388894
rect 423586 388658 423822 388894
rect 423266 388338 423502 388574
rect 423586 388338 423822 388574
rect 185410 381218 185646 381454
rect 185410 380898 185646 381134
rect 216130 381218 216366 381454
rect 216130 380898 216366 381134
rect 246850 381218 247086 381454
rect 246850 380898 247086 381134
rect 277570 381218 277806 381454
rect 277570 380898 277806 381134
rect 308290 381218 308526 381454
rect 308290 380898 308526 381134
rect 339010 381218 339246 381454
rect 339010 380898 339246 381134
rect 369730 381218 369966 381454
rect 369730 380898 369966 381134
rect 400450 381218 400686 381454
rect 400450 380898 400686 381134
rect 156986 374378 157222 374614
rect 157306 374378 157542 374614
rect 156986 374058 157222 374294
rect 157306 374058 157542 374294
rect 170050 363218 170286 363454
rect 170050 362898 170286 363134
rect 200770 363218 201006 363454
rect 200770 362898 201006 363134
rect 231490 363218 231726 363454
rect 231490 362898 231726 363134
rect 262210 363218 262446 363454
rect 262210 362898 262446 363134
rect 292930 363218 293166 363454
rect 292930 362898 293166 363134
rect 323650 363218 323886 363454
rect 323650 362898 323886 363134
rect 354370 363218 354606 363454
rect 354370 362898 354606 363134
rect 385090 363218 385326 363454
rect 385090 362898 385326 363134
rect 415810 363218 416046 363454
rect 415810 362898 416046 363134
rect 423266 352658 423502 352894
rect 423586 352658 423822 352894
rect 423266 352338 423502 352574
rect 423586 352338 423822 352574
rect 185410 345218 185646 345454
rect 185410 344898 185646 345134
rect 216130 345218 216366 345454
rect 216130 344898 216366 345134
rect 246850 345218 247086 345454
rect 246850 344898 247086 345134
rect 277570 345218 277806 345454
rect 277570 344898 277806 345134
rect 308290 345218 308526 345454
rect 308290 344898 308526 345134
rect 339010 345218 339246 345454
rect 339010 344898 339246 345134
rect 369730 345218 369966 345454
rect 369730 344898 369966 345134
rect 400450 345218 400686 345454
rect 400450 344898 400686 345134
rect 156986 338378 157222 338614
rect 157306 338378 157542 338614
rect 156986 338058 157222 338294
rect 157306 338058 157542 338294
rect 170050 327218 170286 327454
rect 170050 326898 170286 327134
rect 200770 327218 201006 327454
rect 200770 326898 201006 327134
rect 231490 327218 231726 327454
rect 231490 326898 231726 327134
rect 262210 327218 262446 327454
rect 262210 326898 262446 327134
rect 292930 327218 293166 327454
rect 292930 326898 293166 327134
rect 323650 327218 323886 327454
rect 323650 326898 323886 327134
rect 354370 327218 354606 327454
rect 354370 326898 354606 327134
rect 385090 327218 385326 327454
rect 385090 326898 385326 327134
rect 415810 327218 416046 327454
rect 415810 326898 416046 327134
rect 423266 316658 423502 316894
rect 423586 316658 423822 316894
rect 423266 316338 423502 316574
rect 423586 316338 423822 316574
rect 185410 309218 185646 309454
rect 185410 308898 185646 309134
rect 216130 309218 216366 309454
rect 216130 308898 216366 309134
rect 246850 309218 247086 309454
rect 246850 308898 247086 309134
rect 277570 309218 277806 309454
rect 277570 308898 277806 309134
rect 308290 309218 308526 309454
rect 308290 308898 308526 309134
rect 339010 309218 339246 309454
rect 339010 308898 339246 309134
rect 369730 309218 369966 309454
rect 369730 308898 369966 309134
rect 400450 309218 400686 309454
rect 400450 308898 400686 309134
rect 156986 302378 157222 302614
rect 157306 302378 157542 302614
rect 156986 302058 157222 302294
rect 157306 302058 157542 302294
rect 170050 291218 170286 291454
rect 170050 290898 170286 291134
rect 200770 291218 201006 291454
rect 200770 290898 201006 291134
rect 231490 291218 231726 291454
rect 231490 290898 231726 291134
rect 262210 291218 262446 291454
rect 262210 290898 262446 291134
rect 292930 291218 293166 291454
rect 292930 290898 293166 291134
rect 323650 291218 323886 291454
rect 323650 290898 323886 291134
rect 354370 291218 354606 291454
rect 354370 290898 354606 291134
rect 385090 291218 385326 291454
rect 385090 290898 385326 291134
rect 415810 291218 416046 291454
rect 415810 290898 416046 291134
rect 423266 280658 423502 280894
rect 423586 280658 423822 280894
rect 423266 280338 423502 280574
rect 423586 280338 423822 280574
rect 185410 273218 185646 273454
rect 185410 272898 185646 273134
rect 216130 273218 216366 273454
rect 216130 272898 216366 273134
rect 246850 273218 247086 273454
rect 246850 272898 247086 273134
rect 277570 273218 277806 273454
rect 277570 272898 277806 273134
rect 308290 273218 308526 273454
rect 308290 272898 308526 273134
rect 339010 273218 339246 273454
rect 339010 272898 339246 273134
rect 369730 273218 369966 273454
rect 369730 272898 369966 273134
rect 400450 273218 400686 273454
rect 400450 272898 400686 273134
rect 156986 266378 157222 266614
rect 157306 266378 157542 266614
rect 156986 266058 157222 266294
rect 157306 266058 157542 266294
rect 170050 255218 170286 255454
rect 170050 254898 170286 255134
rect 200770 255218 201006 255454
rect 200770 254898 201006 255134
rect 231490 255218 231726 255454
rect 231490 254898 231726 255134
rect 262210 255218 262446 255454
rect 262210 254898 262446 255134
rect 292930 255218 293166 255454
rect 292930 254898 293166 255134
rect 323650 255218 323886 255454
rect 323650 254898 323886 255134
rect 354370 255218 354606 255454
rect 354370 254898 354606 255134
rect 385090 255218 385326 255454
rect 385090 254898 385326 255134
rect 415810 255218 416046 255454
rect 415810 254898 416046 255134
rect 423266 244658 423502 244894
rect 423586 244658 423822 244894
rect 423266 244338 423502 244574
rect 423586 244338 423822 244574
rect 185410 237218 185646 237454
rect 185410 236898 185646 237134
rect 216130 237218 216366 237454
rect 216130 236898 216366 237134
rect 246850 237218 247086 237454
rect 246850 236898 247086 237134
rect 277570 237218 277806 237454
rect 277570 236898 277806 237134
rect 308290 237218 308526 237454
rect 308290 236898 308526 237134
rect 339010 237218 339246 237454
rect 339010 236898 339246 237134
rect 369730 237218 369966 237454
rect 369730 236898 369966 237134
rect 400450 237218 400686 237454
rect 400450 236898 400686 237134
rect 156986 230378 157222 230614
rect 157306 230378 157542 230614
rect 156986 230058 157222 230294
rect 157306 230058 157542 230294
rect 170050 219218 170286 219454
rect 170050 218898 170286 219134
rect 200770 219218 201006 219454
rect 200770 218898 201006 219134
rect 231490 219218 231726 219454
rect 231490 218898 231726 219134
rect 262210 219218 262446 219454
rect 262210 218898 262446 219134
rect 292930 219218 293166 219454
rect 292930 218898 293166 219134
rect 323650 219218 323886 219454
rect 323650 218898 323886 219134
rect 354370 219218 354606 219454
rect 354370 218898 354606 219134
rect 385090 219218 385326 219454
rect 385090 218898 385326 219134
rect 415810 219218 416046 219454
rect 415810 218898 416046 219134
rect 423266 208658 423502 208894
rect 423586 208658 423822 208894
rect 423266 208338 423502 208574
rect 423586 208338 423822 208574
rect 156986 194378 157222 194614
rect 157306 194378 157542 194614
rect 156986 194058 157222 194294
rect 157306 194058 157542 194294
rect 156986 158378 157222 158614
rect 157306 158378 157542 158614
rect 156986 158058 157222 158294
rect 157306 158058 157542 158294
rect 156986 122378 157222 122614
rect 157306 122378 157542 122614
rect 156986 122058 157222 122294
rect 157306 122058 157542 122294
rect 156986 86378 157222 86614
rect 157306 86378 157542 86614
rect 156986 86058 157222 86294
rect 157306 86058 157542 86294
rect 156986 50378 157222 50614
rect 157306 50378 157542 50614
rect 156986 50058 157222 50294
rect 157306 50058 157542 50294
rect 156986 14378 157222 14614
rect 157306 14378 157542 14614
rect 156986 14058 157222 14294
rect 157306 14058 157542 14294
rect 138986 -7302 139222 -7066
rect 139306 -7302 139542 -7066
rect 138986 -7622 139222 -7386
rect 139306 -7622 139542 -7386
rect 163826 165218 164062 165454
rect 164146 165218 164382 165454
rect 163826 164898 164062 165134
rect 164146 164898 164382 165134
rect 163826 129218 164062 129454
rect 164146 129218 164382 129454
rect 163826 128898 164062 129134
rect 164146 128898 164382 129134
rect 163826 93218 164062 93454
rect 164146 93218 164382 93454
rect 163826 92898 164062 93134
rect 164146 92898 164382 93134
rect 163826 57218 164062 57454
rect 164146 57218 164382 57454
rect 163826 56898 164062 57134
rect 164146 56898 164382 57134
rect 163826 21218 164062 21454
rect 164146 21218 164382 21454
rect 163826 20898 164062 21134
rect 164146 20898 164382 21134
rect 163826 -1542 164062 -1306
rect 164146 -1542 164382 -1306
rect 163826 -1862 164062 -1626
rect 164146 -1862 164382 -1626
rect 167546 168938 167782 169174
rect 167866 168938 168102 169174
rect 167546 168618 167782 168854
rect 167866 168618 168102 168854
rect 167546 132938 167782 133174
rect 167866 132938 168102 133174
rect 167546 132618 167782 132854
rect 167866 132618 168102 132854
rect 167546 96938 167782 97174
rect 167866 96938 168102 97174
rect 167546 96618 167782 96854
rect 167866 96618 168102 96854
rect 167546 60938 167782 61174
rect 167866 60938 168102 61174
rect 167546 60618 167782 60854
rect 167866 60618 168102 60854
rect 167546 24938 167782 25174
rect 167866 24938 168102 25174
rect 167546 24618 167782 24854
rect 167866 24618 168102 24854
rect 167546 -3462 167782 -3226
rect 167866 -3462 168102 -3226
rect 167546 -3782 167782 -3546
rect 167866 -3782 168102 -3546
rect 171266 172658 171502 172894
rect 171586 172658 171822 172894
rect 171266 172338 171502 172574
rect 171586 172338 171822 172574
rect 171266 136658 171502 136894
rect 171586 136658 171822 136894
rect 171266 136338 171502 136574
rect 171586 136338 171822 136574
rect 171266 100658 171502 100894
rect 171586 100658 171822 100894
rect 171266 100338 171502 100574
rect 171586 100338 171822 100574
rect 171266 64658 171502 64894
rect 171586 64658 171822 64894
rect 171266 64338 171502 64574
rect 171586 64338 171822 64574
rect 171266 28658 171502 28894
rect 171586 28658 171822 28894
rect 171266 28338 171502 28574
rect 171586 28338 171822 28574
rect 171266 -5382 171502 -5146
rect 171586 -5382 171822 -5146
rect 171266 -5702 171502 -5466
rect 171586 -5702 171822 -5466
rect 174986 176378 175222 176614
rect 175306 176378 175542 176614
rect 174986 176058 175222 176294
rect 175306 176058 175542 176294
rect 174986 140378 175222 140614
rect 175306 140378 175542 140614
rect 174986 140058 175222 140294
rect 175306 140058 175542 140294
rect 174986 104378 175222 104614
rect 175306 104378 175542 104614
rect 174986 104058 175222 104294
rect 175306 104058 175542 104294
rect 174986 68378 175222 68614
rect 175306 68378 175542 68614
rect 174986 68058 175222 68294
rect 175306 68058 175542 68294
rect 174986 32378 175222 32614
rect 175306 32378 175542 32614
rect 174986 32058 175222 32294
rect 175306 32058 175542 32294
rect 156986 -6342 157222 -6106
rect 157306 -6342 157542 -6106
rect 156986 -6662 157222 -6426
rect 157306 -6662 157542 -6426
rect 181826 183218 182062 183454
rect 182146 183218 182382 183454
rect 181826 182898 182062 183134
rect 182146 182898 182382 183134
rect 181826 147218 182062 147454
rect 182146 147218 182382 147454
rect 181826 146898 182062 147134
rect 182146 146898 182382 147134
rect 181826 111218 182062 111454
rect 182146 111218 182382 111454
rect 181826 110898 182062 111134
rect 182146 110898 182382 111134
rect 181826 75218 182062 75454
rect 182146 75218 182382 75454
rect 181826 74898 182062 75134
rect 182146 74898 182382 75134
rect 181826 39218 182062 39454
rect 182146 39218 182382 39454
rect 181826 38898 182062 39134
rect 182146 38898 182382 39134
rect 181826 3218 182062 3454
rect 182146 3218 182382 3454
rect 181826 2898 182062 3134
rect 182146 2898 182382 3134
rect 181826 -582 182062 -346
rect 182146 -582 182382 -346
rect 181826 -902 182062 -666
rect 182146 -902 182382 -666
rect 185546 186938 185782 187174
rect 185866 186938 186102 187174
rect 185546 186618 185782 186854
rect 185866 186618 186102 186854
rect 185546 150938 185782 151174
rect 185866 150938 186102 151174
rect 185546 150618 185782 150854
rect 185866 150618 186102 150854
rect 185546 114938 185782 115174
rect 185866 114938 186102 115174
rect 185546 114618 185782 114854
rect 185866 114618 186102 114854
rect 185546 78938 185782 79174
rect 185866 78938 186102 79174
rect 185546 78618 185782 78854
rect 185866 78618 186102 78854
rect 185546 42938 185782 43174
rect 185866 42938 186102 43174
rect 185546 42618 185782 42854
rect 185866 42618 186102 42854
rect 185546 6938 185782 7174
rect 185866 6938 186102 7174
rect 185546 6618 185782 6854
rect 185866 6618 186102 6854
rect 185546 -2502 185782 -2266
rect 185866 -2502 186102 -2266
rect 185546 -2822 185782 -2586
rect 185866 -2822 186102 -2586
rect 189266 190658 189502 190894
rect 189586 190658 189822 190894
rect 189266 190338 189502 190574
rect 189586 190338 189822 190574
rect 189266 154658 189502 154894
rect 189586 154658 189822 154894
rect 189266 154338 189502 154574
rect 189586 154338 189822 154574
rect 189266 118658 189502 118894
rect 189586 118658 189822 118894
rect 189266 118338 189502 118574
rect 189586 118338 189822 118574
rect 189266 82658 189502 82894
rect 189586 82658 189822 82894
rect 189266 82338 189502 82574
rect 189586 82338 189822 82574
rect 189266 46658 189502 46894
rect 189586 46658 189822 46894
rect 189266 46338 189502 46574
rect 189586 46338 189822 46574
rect 189266 10658 189502 10894
rect 189586 10658 189822 10894
rect 189266 10338 189502 10574
rect 189586 10338 189822 10574
rect 189266 -4422 189502 -4186
rect 189586 -4422 189822 -4186
rect 189266 -4742 189502 -4506
rect 189586 -4742 189822 -4506
rect 192986 194378 193222 194614
rect 193306 194378 193542 194614
rect 192986 194058 193222 194294
rect 193306 194058 193542 194294
rect 192986 158378 193222 158614
rect 193306 158378 193542 158614
rect 192986 158058 193222 158294
rect 193306 158058 193542 158294
rect 192986 122378 193222 122614
rect 193306 122378 193542 122614
rect 192986 122058 193222 122294
rect 193306 122058 193542 122294
rect 192986 86378 193222 86614
rect 193306 86378 193542 86614
rect 192986 86058 193222 86294
rect 193306 86058 193542 86294
rect 192986 50378 193222 50614
rect 193306 50378 193542 50614
rect 192986 50058 193222 50294
rect 193306 50058 193542 50294
rect 192986 14378 193222 14614
rect 193306 14378 193542 14614
rect 192986 14058 193222 14294
rect 193306 14058 193542 14294
rect 174986 -7302 175222 -7066
rect 175306 -7302 175542 -7066
rect 174986 -7622 175222 -7386
rect 175306 -7622 175542 -7386
rect 199826 165218 200062 165454
rect 200146 165218 200382 165454
rect 199826 164898 200062 165134
rect 200146 164898 200382 165134
rect 199826 129218 200062 129454
rect 200146 129218 200382 129454
rect 199826 128898 200062 129134
rect 200146 128898 200382 129134
rect 199826 93218 200062 93454
rect 200146 93218 200382 93454
rect 199826 92898 200062 93134
rect 200146 92898 200382 93134
rect 199826 57218 200062 57454
rect 200146 57218 200382 57454
rect 199826 56898 200062 57134
rect 200146 56898 200382 57134
rect 199826 21218 200062 21454
rect 200146 21218 200382 21454
rect 199826 20898 200062 21134
rect 200146 20898 200382 21134
rect 199826 -1542 200062 -1306
rect 200146 -1542 200382 -1306
rect 199826 -1862 200062 -1626
rect 200146 -1862 200382 -1626
rect 203546 168938 203782 169174
rect 203866 168938 204102 169174
rect 203546 168618 203782 168854
rect 203866 168618 204102 168854
rect 203546 132938 203782 133174
rect 203866 132938 204102 133174
rect 203546 132618 203782 132854
rect 203866 132618 204102 132854
rect 203546 96938 203782 97174
rect 203866 96938 204102 97174
rect 203546 96618 203782 96854
rect 203866 96618 204102 96854
rect 203546 60938 203782 61174
rect 203866 60938 204102 61174
rect 203546 60618 203782 60854
rect 203866 60618 204102 60854
rect 203546 24938 203782 25174
rect 203866 24938 204102 25174
rect 203546 24618 203782 24854
rect 203866 24618 204102 24854
rect 203546 -3462 203782 -3226
rect 203866 -3462 204102 -3226
rect 203546 -3782 203782 -3546
rect 203866 -3782 204102 -3546
rect 207266 172658 207502 172894
rect 207586 172658 207822 172894
rect 207266 172338 207502 172574
rect 207586 172338 207822 172574
rect 207266 136658 207502 136894
rect 207586 136658 207822 136894
rect 207266 136338 207502 136574
rect 207586 136338 207822 136574
rect 207266 100658 207502 100894
rect 207586 100658 207822 100894
rect 207266 100338 207502 100574
rect 207586 100338 207822 100574
rect 207266 64658 207502 64894
rect 207586 64658 207822 64894
rect 207266 64338 207502 64574
rect 207586 64338 207822 64574
rect 207266 28658 207502 28894
rect 207586 28658 207822 28894
rect 207266 28338 207502 28574
rect 207586 28338 207822 28574
rect 207266 -5382 207502 -5146
rect 207586 -5382 207822 -5146
rect 207266 -5702 207502 -5466
rect 207586 -5702 207822 -5466
rect 210986 176378 211222 176614
rect 211306 176378 211542 176614
rect 210986 176058 211222 176294
rect 211306 176058 211542 176294
rect 210986 140378 211222 140614
rect 211306 140378 211542 140614
rect 210986 140058 211222 140294
rect 211306 140058 211542 140294
rect 210986 104378 211222 104614
rect 211306 104378 211542 104614
rect 210986 104058 211222 104294
rect 211306 104058 211542 104294
rect 210986 68378 211222 68614
rect 211306 68378 211542 68614
rect 210986 68058 211222 68294
rect 211306 68058 211542 68294
rect 210986 32378 211222 32614
rect 211306 32378 211542 32614
rect 210986 32058 211222 32294
rect 211306 32058 211542 32294
rect 192986 -6342 193222 -6106
rect 193306 -6342 193542 -6106
rect 192986 -6662 193222 -6426
rect 193306 -6662 193542 -6426
rect 217826 183218 218062 183454
rect 218146 183218 218382 183454
rect 217826 182898 218062 183134
rect 218146 182898 218382 183134
rect 217826 147218 218062 147454
rect 218146 147218 218382 147454
rect 217826 146898 218062 147134
rect 218146 146898 218382 147134
rect 217826 111218 218062 111454
rect 218146 111218 218382 111454
rect 217826 110898 218062 111134
rect 218146 110898 218382 111134
rect 217826 75218 218062 75454
rect 218146 75218 218382 75454
rect 217826 74898 218062 75134
rect 218146 74898 218382 75134
rect 217826 39218 218062 39454
rect 218146 39218 218382 39454
rect 217826 38898 218062 39134
rect 218146 38898 218382 39134
rect 217826 3218 218062 3454
rect 218146 3218 218382 3454
rect 217826 2898 218062 3134
rect 218146 2898 218382 3134
rect 217826 -582 218062 -346
rect 218146 -582 218382 -346
rect 217826 -902 218062 -666
rect 218146 -902 218382 -666
rect 221546 186938 221782 187174
rect 221866 186938 222102 187174
rect 221546 186618 221782 186854
rect 221866 186618 222102 186854
rect 221546 150938 221782 151174
rect 221866 150938 222102 151174
rect 221546 150618 221782 150854
rect 221866 150618 222102 150854
rect 221546 114938 221782 115174
rect 221866 114938 222102 115174
rect 221546 114618 221782 114854
rect 221866 114618 222102 114854
rect 221546 78938 221782 79174
rect 221866 78938 222102 79174
rect 221546 78618 221782 78854
rect 221866 78618 222102 78854
rect 221546 42938 221782 43174
rect 221866 42938 222102 43174
rect 221546 42618 221782 42854
rect 221866 42618 222102 42854
rect 221546 6938 221782 7174
rect 221866 6938 222102 7174
rect 221546 6618 221782 6854
rect 221866 6618 222102 6854
rect 221546 -2502 221782 -2266
rect 221866 -2502 222102 -2266
rect 221546 -2822 221782 -2586
rect 221866 -2822 222102 -2586
rect 225266 190658 225502 190894
rect 225586 190658 225822 190894
rect 225266 190338 225502 190574
rect 225586 190338 225822 190574
rect 225266 154658 225502 154894
rect 225586 154658 225822 154894
rect 225266 154338 225502 154574
rect 225586 154338 225822 154574
rect 225266 118658 225502 118894
rect 225586 118658 225822 118894
rect 225266 118338 225502 118574
rect 225586 118338 225822 118574
rect 225266 82658 225502 82894
rect 225586 82658 225822 82894
rect 225266 82338 225502 82574
rect 225586 82338 225822 82574
rect 225266 46658 225502 46894
rect 225586 46658 225822 46894
rect 225266 46338 225502 46574
rect 225586 46338 225822 46574
rect 225266 10658 225502 10894
rect 225586 10658 225822 10894
rect 225266 10338 225502 10574
rect 225586 10338 225822 10574
rect 225266 -4422 225502 -4186
rect 225586 -4422 225822 -4186
rect 225266 -4742 225502 -4506
rect 225586 -4742 225822 -4506
rect 228986 194378 229222 194614
rect 229306 194378 229542 194614
rect 228986 194058 229222 194294
rect 229306 194058 229542 194294
rect 228986 158378 229222 158614
rect 229306 158378 229542 158614
rect 228986 158058 229222 158294
rect 229306 158058 229542 158294
rect 228986 122378 229222 122614
rect 229306 122378 229542 122614
rect 228986 122058 229222 122294
rect 229306 122058 229542 122294
rect 228986 86378 229222 86614
rect 229306 86378 229542 86614
rect 228986 86058 229222 86294
rect 229306 86058 229542 86294
rect 228986 50378 229222 50614
rect 229306 50378 229542 50614
rect 228986 50058 229222 50294
rect 229306 50058 229542 50294
rect 228986 14378 229222 14614
rect 229306 14378 229542 14614
rect 228986 14058 229222 14294
rect 229306 14058 229542 14294
rect 210986 -7302 211222 -7066
rect 211306 -7302 211542 -7066
rect 210986 -7622 211222 -7386
rect 211306 -7622 211542 -7386
rect 235826 165218 236062 165454
rect 236146 165218 236382 165454
rect 235826 164898 236062 165134
rect 236146 164898 236382 165134
rect 235826 129218 236062 129454
rect 236146 129218 236382 129454
rect 235826 128898 236062 129134
rect 236146 128898 236382 129134
rect 235826 93218 236062 93454
rect 236146 93218 236382 93454
rect 235826 92898 236062 93134
rect 236146 92898 236382 93134
rect 235826 57218 236062 57454
rect 236146 57218 236382 57454
rect 235826 56898 236062 57134
rect 236146 56898 236382 57134
rect 235826 21218 236062 21454
rect 236146 21218 236382 21454
rect 235826 20898 236062 21134
rect 236146 20898 236382 21134
rect 235826 -1542 236062 -1306
rect 236146 -1542 236382 -1306
rect 235826 -1862 236062 -1626
rect 236146 -1862 236382 -1626
rect 239546 168938 239782 169174
rect 239866 168938 240102 169174
rect 239546 168618 239782 168854
rect 239866 168618 240102 168854
rect 239546 132938 239782 133174
rect 239866 132938 240102 133174
rect 239546 132618 239782 132854
rect 239866 132618 240102 132854
rect 239546 96938 239782 97174
rect 239866 96938 240102 97174
rect 239546 96618 239782 96854
rect 239866 96618 240102 96854
rect 239546 60938 239782 61174
rect 239866 60938 240102 61174
rect 239546 60618 239782 60854
rect 239866 60618 240102 60854
rect 239546 24938 239782 25174
rect 239866 24938 240102 25174
rect 239546 24618 239782 24854
rect 239866 24618 240102 24854
rect 239546 -3462 239782 -3226
rect 239866 -3462 240102 -3226
rect 239546 -3782 239782 -3546
rect 239866 -3782 240102 -3546
rect 243266 172658 243502 172894
rect 243586 172658 243822 172894
rect 243266 172338 243502 172574
rect 243586 172338 243822 172574
rect 243266 136658 243502 136894
rect 243586 136658 243822 136894
rect 243266 136338 243502 136574
rect 243586 136338 243822 136574
rect 243266 100658 243502 100894
rect 243586 100658 243822 100894
rect 243266 100338 243502 100574
rect 243586 100338 243822 100574
rect 243266 64658 243502 64894
rect 243586 64658 243822 64894
rect 243266 64338 243502 64574
rect 243586 64338 243822 64574
rect 243266 28658 243502 28894
rect 243586 28658 243822 28894
rect 243266 28338 243502 28574
rect 243586 28338 243822 28574
rect 243266 -5382 243502 -5146
rect 243586 -5382 243822 -5146
rect 243266 -5702 243502 -5466
rect 243586 -5702 243822 -5466
rect 246986 176378 247222 176614
rect 247306 176378 247542 176614
rect 246986 176058 247222 176294
rect 247306 176058 247542 176294
rect 246986 140378 247222 140614
rect 247306 140378 247542 140614
rect 246986 140058 247222 140294
rect 247306 140058 247542 140294
rect 246986 104378 247222 104614
rect 247306 104378 247542 104614
rect 246986 104058 247222 104294
rect 247306 104058 247542 104294
rect 246986 68378 247222 68614
rect 247306 68378 247542 68614
rect 246986 68058 247222 68294
rect 247306 68058 247542 68294
rect 246986 32378 247222 32614
rect 247306 32378 247542 32614
rect 246986 32058 247222 32294
rect 247306 32058 247542 32294
rect 228986 -6342 229222 -6106
rect 229306 -6342 229542 -6106
rect 228986 -6662 229222 -6426
rect 229306 -6662 229542 -6426
rect 253826 183218 254062 183454
rect 254146 183218 254382 183454
rect 253826 182898 254062 183134
rect 254146 182898 254382 183134
rect 253826 147218 254062 147454
rect 254146 147218 254382 147454
rect 253826 146898 254062 147134
rect 254146 146898 254382 147134
rect 253826 111218 254062 111454
rect 254146 111218 254382 111454
rect 253826 110898 254062 111134
rect 254146 110898 254382 111134
rect 253826 75218 254062 75454
rect 254146 75218 254382 75454
rect 253826 74898 254062 75134
rect 254146 74898 254382 75134
rect 253826 39218 254062 39454
rect 254146 39218 254382 39454
rect 253826 38898 254062 39134
rect 254146 38898 254382 39134
rect 253826 3218 254062 3454
rect 254146 3218 254382 3454
rect 253826 2898 254062 3134
rect 254146 2898 254382 3134
rect 253826 -582 254062 -346
rect 254146 -582 254382 -346
rect 253826 -902 254062 -666
rect 254146 -902 254382 -666
rect 257546 186938 257782 187174
rect 257866 186938 258102 187174
rect 257546 186618 257782 186854
rect 257866 186618 258102 186854
rect 257546 150938 257782 151174
rect 257866 150938 258102 151174
rect 257546 150618 257782 150854
rect 257866 150618 258102 150854
rect 257546 114938 257782 115174
rect 257866 114938 258102 115174
rect 257546 114618 257782 114854
rect 257866 114618 258102 114854
rect 257546 78938 257782 79174
rect 257866 78938 258102 79174
rect 257546 78618 257782 78854
rect 257866 78618 258102 78854
rect 257546 42938 257782 43174
rect 257866 42938 258102 43174
rect 257546 42618 257782 42854
rect 257866 42618 258102 42854
rect 257546 6938 257782 7174
rect 257866 6938 258102 7174
rect 257546 6618 257782 6854
rect 257866 6618 258102 6854
rect 257546 -2502 257782 -2266
rect 257866 -2502 258102 -2266
rect 257546 -2822 257782 -2586
rect 257866 -2822 258102 -2586
rect 261266 190658 261502 190894
rect 261586 190658 261822 190894
rect 261266 190338 261502 190574
rect 261586 190338 261822 190574
rect 261266 154658 261502 154894
rect 261586 154658 261822 154894
rect 261266 154338 261502 154574
rect 261586 154338 261822 154574
rect 261266 118658 261502 118894
rect 261586 118658 261822 118894
rect 261266 118338 261502 118574
rect 261586 118338 261822 118574
rect 261266 82658 261502 82894
rect 261586 82658 261822 82894
rect 261266 82338 261502 82574
rect 261586 82338 261822 82574
rect 261266 46658 261502 46894
rect 261586 46658 261822 46894
rect 261266 46338 261502 46574
rect 261586 46338 261822 46574
rect 261266 10658 261502 10894
rect 261586 10658 261822 10894
rect 261266 10338 261502 10574
rect 261586 10338 261822 10574
rect 261266 -4422 261502 -4186
rect 261586 -4422 261822 -4186
rect 261266 -4742 261502 -4506
rect 261586 -4742 261822 -4506
rect 264986 194378 265222 194614
rect 265306 194378 265542 194614
rect 264986 194058 265222 194294
rect 265306 194058 265542 194294
rect 264986 158378 265222 158614
rect 265306 158378 265542 158614
rect 264986 158058 265222 158294
rect 265306 158058 265542 158294
rect 264986 122378 265222 122614
rect 265306 122378 265542 122614
rect 264986 122058 265222 122294
rect 265306 122058 265542 122294
rect 264986 86378 265222 86614
rect 265306 86378 265542 86614
rect 264986 86058 265222 86294
rect 265306 86058 265542 86294
rect 264986 50378 265222 50614
rect 265306 50378 265542 50614
rect 264986 50058 265222 50294
rect 265306 50058 265542 50294
rect 264986 14378 265222 14614
rect 265306 14378 265542 14614
rect 264986 14058 265222 14294
rect 265306 14058 265542 14294
rect 246986 -7302 247222 -7066
rect 247306 -7302 247542 -7066
rect 246986 -7622 247222 -7386
rect 247306 -7622 247542 -7386
rect 271826 165218 272062 165454
rect 272146 165218 272382 165454
rect 271826 164898 272062 165134
rect 272146 164898 272382 165134
rect 271826 129218 272062 129454
rect 272146 129218 272382 129454
rect 271826 128898 272062 129134
rect 272146 128898 272382 129134
rect 271826 93218 272062 93454
rect 272146 93218 272382 93454
rect 271826 92898 272062 93134
rect 272146 92898 272382 93134
rect 271826 57218 272062 57454
rect 272146 57218 272382 57454
rect 271826 56898 272062 57134
rect 272146 56898 272382 57134
rect 271826 21218 272062 21454
rect 272146 21218 272382 21454
rect 271826 20898 272062 21134
rect 272146 20898 272382 21134
rect 271826 -1542 272062 -1306
rect 272146 -1542 272382 -1306
rect 271826 -1862 272062 -1626
rect 272146 -1862 272382 -1626
rect 275546 168938 275782 169174
rect 275866 168938 276102 169174
rect 275546 168618 275782 168854
rect 275866 168618 276102 168854
rect 275546 132938 275782 133174
rect 275866 132938 276102 133174
rect 275546 132618 275782 132854
rect 275866 132618 276102 132854
rect 275546 96938 275782 97174
rect 275866 96938 276102 97174
rect 275546 96618 275782 96854
rect 275866 96618 276102 96854
rect 275546 60938 275782 61174
rect 275866 60938 276102 61174
rect 275546 60618 275782 60854
rect 275866 60618 276102 60854
rect 275546 24938 275782 25174
rect 275866 24938 276102 25174
rect 275546 24618 275782 24854
rect 275866 24618 276102 24854
rect 275546 -3462 275782 -3226
rect 275866 -3462 276102 -3226
rect 275546 -3782 275782 -3546
rect 275866 -3782 276102 -3546
rect 279266 172658 279502 172894
rect 279586 172658 279822 172894
rect 279266 172338 279502 172574
rect 279586 172338 279822 172574
rect 279266 136658 279502 136894
rect 279586 136658 279822 136894
rect 279266 136338 279502 136574
rect 279586 136338 279822 136574
rect 279266 100658 279502 100894
rect 279586 100658 279822 100894
rect 279266 100338 279502 100574
rect 279586 100338 279822 100574
rect 279266 64658 279502 64894
rect 279586 64658 279822 64894
rect 279266 64338 279502 64574
rect 279586 64338 279822 64574
rect 279266 28658 279502 28894
rect 279586 28658 279822 28894
rect 279266 28338 279502 28574
rect 279586 28338 279822 28574
rect 279266 -5382 279502 -5146
rect 279586 -5382 279822 -5146
rect 279266 -5702 279502 -5466
rect 279586 -5702 279822 -5466
rect 282986 176378 283222 176614
rect 283306 176378 283542 176614
rect 282986 176058 283222 176294
rect 283306 176058 283542 176294
rect 282986 140378 283222 140614
rect 283306 140378 283542 140614
rect 282986 140058 283222 140294
rect 283306 140058 283542 140294
rect 282986 104378 283222 104614
rect 283306 104378 283542 104614
rect 282986 104058 283222 104294
rect 283306 104058 283542 104294
rect 282986 68378 283222 68614
rect 283306 68378 283542 68614
rect 282986 68058 283222 68294
rect 283306 68058 283542 68294
rect 282986 32378 283222 32614
rect 283306 32378 283542 32614
rect 282986 32058 283222 32294
rect 283306 32058 283542 32294
rect 264986 -6342 265222 -6106
rect 265306 -6342 265542 -6106
rect 264986 -6662 265222 -6426
rect 265306 -6662 265542 -6426
rect 289826 183218 290062 183454
rect 290146 183218 290382 183454
rect 289826 182898 290062 183134
rect 290146 182898 290382 183134
rect 289826 147218 290062 147454
rect 290146 147218 290382 147454
rect 289826 146898 290062 147134
rect 290146 146898 290382 147134
rect 289826 111218 290062 111454
rect 290146 111218 290382 111454
rect 289826 110898 290062 111134
rect 290146 110898 290382 111134
rect 289826 75218 290062 75454
rect 290146 75218 290382 75454
rect 289826 74898 290062 75134
rect 290146 74898 290382 75134
rect 289826 39218 290062 39454
rect 290146 39218 290382 39454
rect 289826 38898 290062 39134
rect 290146 38898 290382 39134
rect 289826 3218 290062 3454
rect 290146 3218 290382 3454
rect 289826 2898 290062 3134
rect 290146 2898 290382 3134
rect 289826 -582 290062 -346
rect 290146 -582 290382 -346
rect 289826 -902 290062 -666
rect 290146 -902 290382 -666
rect 293546 186938 293782 187174
rect 293866 186938 294102 187174
rect 293546 186618 293782 186854
rect 293866 186618 294102 186854
rect 293546 150938 293782 151174
rect 293866 150938 294102 151174
rect 293546 150618 293782 150854
rect 293866 150618 294102 150854
rect 293546 114938 293782 115174
rect 293866 114938 294102 115174
rect 293546 114618 293782 114854
rect 293866 114618 294102 114854
rect 293546 78938 293782 79174
rect 293866 78938 294102 79174
rect 293546 78618 293782 78854
rect 293866 78618 294102 78854
rect 293546 42938 293782 43174
rect 293866 42938 294102 43174
rect 293546 42618 293782 42854
rect 293866 42618 294102 42854
rect 293546 6938 293782 7174
rect 293866 6938 294102 7174
rect 293546 6618 293782 6854
rect 293866 6618 294102 6854
rect 293546 -2502 293782 -2266
rect 293866 -2502 294102 -2266
rect 293546 -2822 293782 -2586
rect 293866 -2822 294102 -2586
rect 297266 190658 297502 190894
rect 297586 190658 297822 190894
rect 297266 190338 297502 190574
rect 297586 190338 297822 190574
rect 297266 154658 297502 154894
rect 297586 154658 297822 154894
rect 297266 154338 297502 154574
rect 297586 154338 297822 154574
rect 297266 118658 297502 118894
rect 297586 118658 297822 118894
rect 297266 118338 297502 118574
rect 297586 118338 297822 118574
rect 297266 82658 297502 82894
rect 297586 82658 297822 82894
rect 297266 82338 297502 82574
rect 297586 82338 297822 82574
rect 297266 46658 297502 46894
rect 297586 46658 297822 46894
rect 297266 46338 297502 46574
rect 297586 46338 297822 46574
rect 297266 10658 297502 10894
rect 297586 10658 297822 10894
rect 297266 10338 297502 10574
rect 297586 10338 297822 10574
rect 297266 -4422 297502 -4186
rect 297586 -4422 297822 -4186
rect 297266 -4742 297502 -4506
rect 297586 -4742 297822 -4506
rect 300986 194378 301222 194614
rect 301306 194378 301542 194614
rect 300986 194058 301222 194294
rect 301306 194058 301542 194294
rect 300986 158378 301222 158614
rect 301306 158378 301542 158614
rect 300986 158058 301222 158294
rect 301306 158058 301542 158294
rect 300986 122378 301222 122614
rect 301306 122378 301542 122614
rect 300986 122058 301222 122294
rect 301306 122058 301542 122294
rect 300986 86378 301222 86614
rect 301306 86378 301542 86614
rect 300986 86058 301222 86294
rect 301306 86058 301542 86294
rect 300986 50378 301222 50614
rect 301306 50378 301542 50614
rect 300986 50058 301222 50294
rect 301306 50058 301542 50294
rect 300986 14378 301222 14614
rect 301306 14378 301542 14614
rect 300986 14058 301222 14294
rect 301306 14058 301542 14294
rect 282986 -7302 283222 -7066
rect 283306 -7302 283542 -7066
rect 282986 -7622 283222 -7386
rect 283306 -7622 283542 -7386
rect 307826 165218 308062 165454
rect 308146 165218 308382 165454
rect 307826 164898 308062 165134
rect 308146 164898 308382 165134
rect 307826 129218 308062 129454
rect 308146 129218 308382 129454
rect 307826 128898 308062 129134
rect 308146 128898 308382 129134
rect 307826 93218 308062 93454
rect 308146 93218 308382 93454
rect 307826 92898 308062 93134
rect 308146 92898 308382 93134
rect 307826 57218 308062 57454
rect 308146 57218 308382 57454
rect 307826 56898 308062 57134
rect 308146 56898 308382 57134
rect 307826 21218 308062 21454
rect 308146 21218 308382 21454
rect 307826 20898 308062 21134
rect 308146 20898 308382 21134
rect 307826 -1542 308062 -1306
rect 308146 -1542 308382 -1306
rect 307826 -1862 308062 -1626
rect 308146 -1862 308382 -1626
rect 311546 168938 311782 169174
rect 311866 168938 312102 169174
rect 311546 168618 311782 168854
rect 311866 168618 312102 168854
rect 311546 132938 311782 133174
rect 311866 132938 312102 133174
rect 311546 132618 311782 132854
rect 311866 132618 312102 132854
rect 311546 96938 311782 97174
rect 311866 96938 312102 97174
rect 311546 96618 311782 96854
rect 311866 96618 312102 96854
rect 311546 60938 311782 61174
rect 311866 60938 312102 61174
rect 311546 60618 311782 60854
rect 311866 60618 312102 60854
rect 311546 24938 311782 25174
rect 311866 24938 312102 25174
rect 311546 24618 311782 24854
rect 311866 24618 312102 24854
rect 311546 -3462 311782 -3226
rect 311866 -3462 312102 -3226
rect 311546 -3782 311782 -3546
rect 311866 -3782 312102 -3546
rect 315266 172658 315502 172894
rect 315586 172658 315822 172894
rect 315266 172338 315502 172574
rect 315586 172338 315822 172574
rect 315266 136658 315502 136894
rect 315586 136658 315822 136894
rect 315266 136338 315502 136574
rect 315586 136338 315822 136574
rect 315266 100658 315502 100894
rect 315586 100658 315822 100894
rect 315266 100338 315502 100574
rect 315586 100338 315822 100574
rect 315266 64658 315502 64894
rect 315586 64658 315822 64894
rect 315266 64338 315502 64574
rect 315586 64338 315822 64574
rect 315266 28658 315502 28894
rect 315586 28658 315822 28894
rect 315266 28338 315502 28574
rect 315586 28338 315822 28574
rect 315266 -5382 315502 -5146
rect 315586 -5382 315822 -5146
rect 315266 -5702 315502 -5466
rect 315586 -5702 315822 -5466
rect 318986 176378 319222 176614
rect 319306 176378 319542 176614
rect 318986 176058 319222 176294
rect 319306 176058 319542 176294
rect 318986 140378 319222 140614
rect 319306 140378 319542 140614
rect 318986 140058 319222 140294
rect 319306 140058 319542 140294
rect 318986 104378 319222 104614
rect 319306 104378 319542 104614
rect 318986 104058 319222 104294
rect 319306 104058 319542 104294
rect 318986 68378 319222 68614
rect 319306 68378 319542 68614
rect 318986 68058 319222 68294
rect 319306 68058 319542 68294
rect 318986 32378 319222 32614
rect 319306 32378 319542 32614
rect 318986 32058 319222 32294
rect 319306 32058 319542 32294
rect 300986 -6342 301222 -6106
rect 301306 -6342 301542 -6106
rect 300986 -6662 301222 -6426
rect 301306 -6662 301542 -6426
rect 325826 183218 326062 183454
rect 326146 183218 326382 183454
rect 325826 182898 326062 183134
rect 326146 182898 326382 183134
rect 325826 147218 326062 147454
rect 326146 147218 326382 147454
rect 325826 146898 326062 147134
rect 326146 146898 326382 147134
rect 325826 111218 326062 111454
rect 326146 111218 326382 111454
rect 325826 110898 326062 111134
rect 326146 110898 326382 111134
rect 325826 75218 326062 75454
rect 326146 75218 326382 75454
rect 325826 74898 326062 75134
rect 326146 74898 326382 75134
rect 325826 39218 326062 39454
rect 326146 39218 326382 39454
rect 325826 38898 326062 39134
rect 326146 38898 326382 39134
rect 325826 3218 326062 3454
rect 326146 3218 326382 3454
rect 325826 2898 326062 3134
rect 326146 2898 326382 3134
rect 325826 -582 326062 -346
rect 326146 -582 326382 -346
rect 325826 -902 326062 -666
rect 326146 -902 326382 -666
rect 329546 186938 329782 187174
rect 329866 186938 330102 187174
rect 329546 186618 329782 186854
rect 329866 186618 330102 186854
rect 329546 150938 329782 151174
rect 329866 150938 330102 151174
rect 329546 150618 329782 150854
rect 329866 150618 330102 150854
rect 329546 114938 329782 115174
rect 329866 114938 330102 115174
rect 329546 114618 329782 114854
rect 329866 114618 330102 114854
rect 329546 78938 329782 79174
rect 329866 78938 330102 79174
rect 329546 78618 329782 78854
rect 329866 78618 330102 78854
rect 329546 42938 329782 43174
rect 329866 42938 330102 43174
rect 329546 42618 329782 42854
rect 329866 42618 330102 42854
rect 329546 6938 329782 7174
rect 329866 6938 330102 7174
rect 329546 6618 329782 6854
rect 329866 6618 330102 6854
rect 329546 -2502 329782 -2266
rect 329866 -2502 330102 -2266
rect 329546 -2822 329782 -2586
rect 329866 -2822 330102 -2586
rect 333266 190658 333502 190894
rect 333586 190658 333822 190894
rect 333266 190338 333502 190574
rect 333586 190338 333822 190574
rect 333266 154658 333502 154894
rect 333586 154658 333822 154894
rect 333266 154338 333502 154574
rect 333586 154338 333822 154574
rect 333266 118658 333502 118894
rect 333586 118658 333822 118894
rect 333266 118338 333502 118574
rect 333586 118338 333822 118574
rect 333266 82658 333502 82894
rect 333586 82658 333822 82894
rect 333266 82338 333502 82574
rect 333586 82338 333822 82574
rect 333266 46658 333502 46894
rect 333586 46658 333822 46894
rect 333266 46338 333502 46574
rect 333586 46338 333822 46574
rect 333266 10658 333502 10894
rect 333586 10658 333822 10894
rect 333266 10338 333502 10574
rect 333586 10338 333822 10574
rect 333266 -4422 333502 -4186
rect 333586 -4422 333822 -4186
rect 333266 -4742 333502 -4506
rect 333586 -4742 333822 -4506
rect 336986 194378 337222 194614
rect 337306 194378 337542 194614
rect 336986 194058 337222 194294
rect 337306 194058 337542 194294
rect 336986 158378 337222 158614
rect 337306 158378 337542 158614
rect 336986 158058 337222 158294
rect 337306 158058 337542 158294
rect 336986 122378 337222 122614
rect 337306 122378 337542 122614
rect 336986 122058 337222 122294
rect 337306 122058 337542 122294
rect 336986 86378 337222 86614
rect 337306 86378 337542 86614
rect 336986 86058 337222 86294
rect 337306 86058 337542 86294
rect 336986 50378 337222 50614
rect 337306 50378 337542 50614
rect 336986 50058 337222 50294
rect 337306 50058 337542 50294
rect 336986 14378 337222 14614
rect 337306 14378 337542 14614
rect 336986 14058 337222 14294
rect 337306 14058 337542 14294
rect 318986 -7302 319222 -7066
rect 319306 -7302 319542 -7066
rect 318986 -7622 319222 -7386
rect 319306 -7622 319542 -7386
rect 343826 165218 344062 165454
rect 344146 165218 344382 165454
rect 343826 164898 344062 165134
rect 344146 164898 344382 165134
rect 343826 129218 344062 129454
rect 344146 129218 344382 129454
rect 343826 128898 344062 129134
rect 344146 128898 344382 129134
rect 343826 93218 344062 93454
rect 344146 93218 344382 93454
rect 343826 92898 344062 93134
rect 344146 92898 344382 93134
rect 343826 57218 344062 57454
rect 344146 57218 344382 57454
rect 343826 56898 344062 57134
rect 344146 56898 344382 57134
rect 343826 21218 344062 21454
rect 344146 21218 344382 21454
rect 343826 20898 344062 21134
rect 344146 20898 344382 21134
rect 343826 -1542 344062 -1306
rect 344146 -1542 344382 -1306
rect 343826 -1862 344062 -1626
rect 344146 -1862 344382 -1626
rect 347546 168938 347782 169174
rect 347866 168938 348102 169174
rect 347546 168618 347782 168854
rect 347866 168618 348102 168854
rect 347546 132938 347782 133174
rect 347866 132938 348102 133174
rect 347546 132618 347782 132854
rect 347866 132618 348102 132854
rect 347546 96938 347782 97174
rect 347866 96938 348102 97174
rect 347546 96618 347782 96854
rect 347866 96618 348102 96854
rect 347546 60938 347782 61174
rect 347866 60938 348102 61174
rect 347546 60618 347782 60854
rect 347866 60618 348102 60854
rect 347546 24938 347782 25174
rect 347866 24938 348102 25174
rect 347546 24618 347782 24854
rect 347866 24618 348102 24854
rect 347546 -3462 347782 -3226
rect 347866 -3462 348102 -3226
rect 347546 -3782 347782 -3546
rect 347866 -3782 348102 -3546
rect 351266 172658 351502 172894
rect 351586 172658 351822 172894
rect 351266 172338 351502 172574
rect 351586 172338 351822 172574
rect 351266 136658 351502 136894
rect 351586 136658 351822 136894
rect 351266 136338 351502 136574
rect 351586 136338 351822 136574
rect 351266 100658 351502 100894
rect 351586 100658 351822 100894
rect 351266 100338 351502 100574
rect 351586 100338 351822 100574
rect 351266 64658 351502 64894
rect 351586 64658 351822 64894
rect 351266 64338 351502 64574
rect 351586 64338 351822 64574
rect 351266 28658 351502 28894
rect 351586 28658 351822 28894
rect 351266 28338 351502 28574
rect 351586 28338 351822 28574
rect 351266 -5382 351502 -5146
rect 351586 -5382 351822 -5146
rect 351266 -5702 351502 -5466
rect 351586 -5702 351822 -5466
rect 354986 176378 355222 176614
rect 355306 176378 355542 176614
rect 354986 176058 355222 176294
rect 355306 176058 355542 176294
rect 354986 140378 355222 140614
rect 355306 140378 355542 140614
rect 354986 140058 355222 140294
rect 355306 140058 355542 140294
rect 354986 104378 355222 104614
rect 355306 104378 355542 104614
rect 354986 104058 355222 104294
rect 355306 104058 355542 104294
rect 354986 68378 355222 68614
rect 355306 68378 355542 68614
rect 354986 68058 355222 68294
rect 355306 68058 355542 68294
rect 354986 32378 355222 32614
rect 355306 32378 355542 32614
rect 354986 32058 355222 32294
rect 355306 32058 355542 32294
rect 336986 -6342 337222 -6106
rect 337306 -6342 337542 -6106
rect 336986 -6662 337222 -6426
rect 337306 -6662 337542 -6426
rect 361826 183218 362062 183454
rect 362146 183218 362382 183454
rect 361826 182898 362062 183134
rect 362146 182898 362382 183134
rect 361826 147218 362062 147454
rect 362146 147218 362382 147454
rect 361826 146898 362062 147134
rect 362146 146898 362382 147134
rect 361826 111218 362062 111454
rect 362146 111218 362382 111454
rect 361826 110898 362062 111134
rect 362146 110898 362382 111134
rect 361826 75218 362062 75454
rect 362146 75218 362382 75454
rect 361826 74898 362062 75134
rect 362146 74898 362382 75134
rect 361826 39218 362062 39454
rect 362146 39218 362382 39454
rect 361826 38898 362062 39134
rect 362146 38898 362382 39134
rect 361826 3218 362062 3454
rect 362146 3218 362382 3454
rect 361826 2898 362062 3134
rect 362146 2898 362382 3134
rect 361826 -582 362062 -346
rect 362146 -582 362382 -346
rect 361826 -902 362062 -666
rect 362146 -902 362382 -666
rect 365546 186938 365782 187174
rect 365866 186938 366102 187174
rect 365546 186618 365782 186854
rect 365866 186618 366102 186854
rect 365546 150938 365782 151174
rect 365866 150938 366102 151174
rect 365546 150618 365782 150854
rect 365866 150618 366102 150854
rect 365546 114938 365782 115174
rect 365866 114938 366102 115174
rect 365546 114618 365782 114854
rect 365866 114618 366102 114854
rect 365546 78938 365782 79174
rect 365866 78938 366102 79174
rect 365546 78618 365782 78854
rect 365866 78618 366102 78854
rect 365546 42938 365782 43174
rect 365866 42938 366102 43174
rect 365546 42618 365782 42854
rect 365866 42618 366102 42854
rect 365546 6938 365782 7174
rect 365866 6938 366102 7174
rect 365546 6618 365782 6854
rect 365866 6618 366102 6854
rect 365546 -2502 365782 -2266
rect 365866 -2502 366102 -2266
rect 365546 -2822 365782 -2586
rect 365866 -2822 366102 -2586
rect 369266 190658 369502 190894
rect 369586 190658 369822 190894
rect 369266 190338 369502 190574
rect 369586 190338 369822 190574
rect 369266 154658 369502 154894
rect 369586 154658 369822 154894
rect 369266 154338 369502 154574
rect 369586 154338 369822 154574
rect 369266 118658 369502 118894
rect 369586 118658 369822 118894
rect 369266 118338 369502 118574
rect 369586 118338 369822 118574
rect 369266 82658 369502 82894
rect 369586 82658 369822 82894
rect 369266 82338 369502 82574
rect 369586 82338 369822 82574
rect 369266 46658 369502 46894
rect 369586 46658 369822 46894
rect 369266 46338 369502 46574
rect 369586 46338 369822 46574
rect 369266 10658 369502 10894
rect 369586 10658 369822 10894
rect 369266 10338 369502 10574
rect 369586 10338 369822 10574
rect 369266 -4422 369502 -4186
rect 369586 -4422 369822 -4186
rect 369266 -4742 369502 -4506
rect 369586 -4742 369822 -4506
rect 372986 194378 373222 194614
rect 373306 194378 373542 194614
rect 372986 194058 373222 194294
rect 373306 194058 373542 194294
rect 372986 158378 373222 158614
rect 373306 158378 373542 158614
rect 372986 158058 373222 158294
rect 373306 158058 373542 158294
rect 372986 122378 373222 122614
rect 373306 122378 373542 122614
rect 372986 122058 373222 122294
rect 373306 122058 373542 122294
rect 372986 86378 373222 86614
rect 373306 86378 373542 86614
rect 372986 86058 373222 86294
rect 373306 86058 373542 86294
rect 372986 50378 373222 50614
rect 373306 50378 373542 50614
rect 372986 50058 373222 50294
rect 373306 50058 373542 50294
rect 372986 14378 373222 14614
rect 373306 14378 373542 14614
rect 372986 14058 373222 14294
rect 373306 14058 373542 14294
rect 354986 -7302 355222 -7066
rect 355306 -7302 355542 -7066
rect 354986 -7622 355222 -7386
rect 355306 -7622 355542 -7386
rect 379826 165218 380062 165454
rect 380146 165218 380382 165454
rect 379826 164898 380062 165134
rect 380146 164898 380382 165134
rect 379826 129218 380062 129454
rect 380146 129218 380382 129454
rect 379826 128898 380062 129134
rect 380146 128898 380382 129134
rect 379826 93218 380062 93454
rect 380146 93218 380382 93454
rect 379826 92898 380062 93134
rect 380146 92898 380382 93134
rect 379826 57218 380062 57454
rect 380146 57218 380382 57454
rect 379826 56898 380062 57134
rect 380146 56898 380382 57134
rect 379826 21218 380062 21454
rect 380146 21218 380382 21454
rect 379826 20898 380062 21134
rect 380146 20898 380382 21134
rect 379826 -1542 380062 -1306
rect 380146 -1542 380382 -1306
rect 379826 -1862 380062 -1626
rect 380146 -1862 380382 -1626
rect 383546 168938 383782 169174
rect 383866 168938 384102 169174
rect 383546 168618 383782 168854
rect 383866 168618 384102 168854
rect 383546 132938 383782 133174
rect 383866 132938 384102 133174
rect 383546 132618 383782 132854
rect 383866 132618 384102 132854
rect 383546 96938 383782 97174
rect 383866 96938 384102 97174
rect 383546 96618 383782 96854
rect 383866 96618 384102 96854
rect 383546 60938 383782 61174
rect 383866 60938 384102 61174
rect 383546 60618 383782 60854
rect 383866 60618 384102 60854
rect 383546 24938 383782 25174
rect 383866 24938 384102 25174
rect 383546 24618 383782 24854
rect 383866 24618 384102 24854
rect 383546 -3462 383782 -3226
rect 383866 -3462 384102 -3226
rect 383546 -3782 383782 -3546
rect 383866 -3782 384102 -3546
rect 387266 172658 387502 172894
rect 387586 172658 387822 172894
rect 387266 172338 387502 172574
rect 387586 172338 387822 172574
rect 387266 136658 387502 136894
rect 387586 136658 387822 136894
rect 387266 136338 387502 136574
rect 387586 136338 387822 136574
rect 387266 100658 387502 100894
rect 387586 100658 387822 100894
rect 387266 100338 387502 100574
rect 387586 100338 387822 100574
rect 387266 64658 387502 64894
rect 387586 64658 387822 64894
rect 387266 64338 387502 64574
rect 387586 64338 387822 64574
rect 387266 28658 387502 28894
rect 387586 28658 387822 28894
rect 387266 28338 387502 28574
rect 387586 28338 387822 28574
rect 387266 -5382 387502 -5146
rect 387586 -5382 387822 -5146
rect 387266 -5702 387502 -5466
rect 387586 -5702 387822 -5466
rect 390986 176378 391222 176614
rect 391306 176378 391542 176614
rect 390986 176058 391222 176294
rect 391306 176058 391542 176294
rect 390986 140378 391222 140614
rect 391306 140378 391542 140614
rect 390986 140058 391222 140294
rect 391306 140058 391542 140294
rect 390986 104378 391222 104614
rect 391306 104378 391542 104614
rect 390986 104058 391222 104294
rect 391306 104058 391542 104294
rect 390986 68378 391222 68614
rect 391306 68378 391542 68614
rect 390986 68058 391222 68294
rect 391306 68058 391542 68294
rect 390986 32378 391222 32614
rect 391306 32378 391542 32614
rect 390986 32058 391222 32294
rect 391306 32058 391542 32294
rect 372986 -6342 373222 -6106
rect 373306 -6342 373542 -6106
rect 372986 -6662 373222 -6426
rect 373306 -6662 373542 -6426
rect 397826 183218 398062 183454
rect 398146 183218 398382 183454
rect 397826 182898 398062 183134
rect 398146 182898 398382 183134
rect 397826 147218 398062 147454
rect 398146 147218 398382 147454
rect 397826 146898 398062 147134
rect 398146 146898 398382 147134
rect 397826 111218 398062 111454
rect 398146 111218 398382 111454
rect 397826 110898 398062 111134
rect 398146 110898 398382 111134
rect 397826 75218 398062 75454
rect 398146 75218 398382 75454
rect 397826 74898 398062 75134
rect 398146 74898 398382 75134
rect 397826 39218 398062 39454
rect 398146 39218 398382 39454
rect 397826 38898 398062 39134
rect 398146 38898 398382 39134
rect 397826 3218 398062 3454
rect 398146 3218 398382 3454
rect 397826 2898 398062 3134
rect 398146 2898 398382 3134
rect 397826 -582 398062 -346
rect 398146 -582 398382 -346
rect 397826 -902 398062 -666
rect 398146 -902 398382 -666
rect 401546 186938 401782 187174
rect 401866 186938 402102 187174
rect 401546 186618 401782 186854
rect 401866 186618 402102 186854
rect 401546 150938 401782 151174
rect 401866 150938 402102 151174
rect 401546 150618 401782 150854
rect 401866 150618 402102 150854
rect 401546 114938 401782 115174
rect 401866 114938 402102 115174
rect 401546 114618 401782 114854
rect 401866 114618 402102 114854
rect 401546 78938 401782 79174
rect 401866 78938 402102 79174
rect 401546 78618 401782 78854
rect 401866 78618 402102 78854
rect 401546 42938 401782 43174
rect 401866 42938 402102 43174
rect 401546 42618 401782 42854
rect 401866 42618 402102 42854
rect 401546 6938 401782 7174
rect 401866 6938 402102 7174
rect 401546 6618 401782 6854
rect 401866 6618 402102 6854
rect 401546 -2502 401782 -2266
rect 401866 -2502 402102 -2266
rect 401546 -2822 401782 -2586
rect 401866 -2822 402102 -2586
rect 405266 190658 405502 190894
rect 405586 190658 405822 190894
rect 405266 190338 405502 190574
rect 405586 190338 405822 190574
rect 405266 154658 405502 154894
rect 405586 154658 405822 154894
rect 405266 154338 405502 154574
rect 405586 154338 405822 154574
rect 405266 118658 405502 118894
rect 405586 118658 405822 118894
rect 405266 118338 405502 118574
rect 405586 118338 405822 118574
rect 405266 82658 405502 82894
rect 405586 82658 405822 82894
rect 405266 82338 405502 82574
rect 405586 82338 405822 82574
rect 405266 46658 405502 46894
rect 405586 46658 405822 46894
rect 405266 46338 405502 46574
rect 405586 46338 405822 46574
rect 405266 10658 405502 10894
rect 405586 10658 405822 10894
rect 405266 10338 405502 10574
rect 405586 10338 405822 10574
rect 405266 -4422 405502 -4186
rect 405586 -4422 405822 -4186
rect 405266 -4742 405502 -4506
rect 405586 -4742 405822 -4506
rect 408986 194378 409222 194614
rect 409306 194378 409542 194614
rect 408986 194058 409222 194294
rect 409306 194058 409542 194294
rect 408986 158378 409222 158614
rect 409306 158378 409542 158614
rect 408986 158058 409222 158294
rect 409306 158058 409542 158294
rect 408986 122378 409222 122614
rect 409306 122378 409542 122614
rect 408986 122058 409222 122294
rect 409306 122058 409542 122294
rect 408986 86378 409222 86614
rect 409306 86378 409542 86614
rect 408986 86058 409222 86294
rect 409306 86058 409542 86294
rect 408986 50378 409222 50614
rect 409306 50378 409542 50614
rect 408986 50058 409222 50294
rect 409306 50058 409542 50294
rect 408986 14378 409222 14614
rect 409306 14378 409542 14614
rect 408986 14058 409222 14294
rect 409306 14058 409542 14294
rect 390986 -7302 391222 -7066
rect 391306 -7302 391542 -7066
rect 390986 -7622 391222 -7386
rect 391306 -7622 391542 -7386
rect 415826 165218 416062 165454
rect 416146 165218 416382 165454
rect 415826 164898 416062 165134
rect 416146 164898 416382 165134
rect 415826 129218 416062 129454
rect 416146 129218 416382 129454
rect 415826 128898 416062 129134
rect 416146 128898 416382 129134
rect 415826 93218 416062 93454
rect 416146 93218 416382 93454
rect 415826 92898 416062 93134
rect 416146 92898 416382 93134
rect 415826 57218 416062 57454
rect 416146 57218 416382 57454
rect 415826 56898 416062 57134
rect 416146 56898 416382 57134
rect 415826 21218 416062 21454
rect 416146 21218 416382 21454
rect 415826 20898 416062 21134
rect 416146 20898 416382 21134
rect 415826 -1542 416062 -1306
rect 416146 -1542 416382 -1306
rect 415826 -1862 416062 -1626
rect 416146 -1862 416382 -1626
rect 419546 168938 419782 169174
rect 419866 168938 420102 169174
rect 419546 168618 419782 168854
rect 419866 168618 420102 168854
rect 419546 132938 419782 133174
rect 419866 132938 420102 133174
rect 419546 132618 419782 132854
rect 419866 132618 420102 132854
rect 419546 96938 419782 97174
rect 419866 96938 420102 97174
rect 419546 96618 419782 96854
rect 419866 96618 420102 96854
rect 419546 60938 419782 61174
rect 419866 60938 420102 61174
rect 419546 60618 419782 60854
rect 419866 60618 420102 60854
rect 419546 24938 419782 25174
rect 419866 24938 420102 25174
rect 419546 24618 419782 24854
rect 419866 24618 420102 24854
rect 419546 -3462 419782 -3226
rect 419866 -3462 420102 -3226
rect 419546 -3782 419782 -3546
rect 419866 -3782 420102 -3546
rect 423266 172658 423502 172894
rect 423586 172658 423822 172894
rect 423266 172338 423502 172574
rect 423586 172338 423822 172574
rect 423266 136658 423502 136894
rect 423586 136658 423822 136894
rect 423266 136338 423502 136574
rect 423586 136338 423822 136574
rect 423266 100658 423502 100894
rect 423586 100658 423822 100894
rect 423266 100338 423502 100574
rect 423586 100338 423822 100574
rect 423266 64658 423502 64894
rect 423586 64658 423822 64894
rect 423266 64338 423502 64574
rect 423586 64338 423822 64574
rect 423266 28658 423502 28894
rect 423586 28658 423822 28894
rect 423266 28338 423502 28574
rect 423586 28338 423822 28574
rect 423266 -5382 423502 -5146
rect 423586 -5382 423822 -5146
rect 423266 -5702 423502 -5466
rect 423586 -5702 423822 -5466
rect 444986 710362 445222 710598
rect 445306 710362 445542 710598
rect 444986 710042 445222 710278
rect 445306 710042 445542 710278
rect 441266 708442 441502 708678
rect 441586 708442 441822 708678
rect 441266 708122 441502 708358
rect 441586 708122 441822 708358
rect 437546 706522 437782 706758
rect 437866 706522 438102 706758
rect 437546 706202 437782 706438
rect 437866 706202 438102 706438
rect 426986 680378 427222 680614
rect 427306 680378 427542 680614
rect 426986 680058 427222 680294
rect 427306 680058 427542 680294
rect 426986 644378 427222 644614
rect 427306 644378 427542 644614
rect 426986 644058 427222 644294
rect 427306 644058 427542 644294
rect 426986 608378 427222 608614
rect 427306 608378 427542 608614
rect 426986 608058 427222 608294
rect 427306 608058 427542 608294
rect 426986 572378 427222 572614
rect 427306 572378 427542 572614
rect 426986 572058 427222 572294
rect 427306 572058 427542 572294
rect 426986 536378 427222 536614
rect 427306 536378 427542 536614
rect 426986 536058 427222 536294
rect 427306 536058 427542 536294
rect 426986 500378 427222 500614
rect 427306 500378 427542 500614
rect 426986 500058 427222 500294
rect 427306 500058 427542 500294
rect 426986 464378 427222 464614
rect 427306 464378 427542 464614
rect 426986 464058 427222 464294
rect 427306 464058 427542 464294
rect 426986 428378 427222 428614
rect 427306 428378 427542 428614
rect 426986 428058 427222 428294
rect 427306 428058 427542 428294
rect 426986 392378 427222 392614
rect 427306 392378 427542 392614
rect 426986 392058 427222 392294
rect 427306 392058 427542 392294
rect 426986 356378 427222 356614
rect 427306 356378 427542 356614
rect 426986 356058 427222 356294
rect 427306 356058 427542 356294
rect 426986 320378 427222 320614
rect 427306 320378 427542 320614
rect 426986 320058 427222 320294
rect 427306 320058 427542 320294
rect 426986 284378 427222 284614
rect 427306 284378 427542 284614
rect 426986 284058 427222 284294
rect 427306 284058 427542 284294
rect 426986 248378 427222 248614
rect 427306 248378 427542 248614
rect 426986 248058 427222 248294
rect 427306 248058 427542 248294
rect 426986 212378 427222 212614
rect 427306 212378 427542 212614
rect 426986 212058 427222 212294
rect 427306 212058 427542 212294
rect 426986 176378 427222 176614
rect 427306 176378 427542 176614
rect 426986 176058 427222 176294
rect 427306 176058 427542 176294
rect 426986 140378 427222 140614
rect 427306 140378 427542 140614
rect 426986 140058 427222 140294
rect 427306 140058 427542 140294
rect 426986 104378 427222 104614
rect 427306 104378 427542 104614
rect 426986 104058 427222 104294
rect 427306 104058 427542 104294
rect 426986 68378 427222 68614
rect 427306 68378 427542 68614
rect 426986 68058 427222 68294
rect 427306 68058 427542 68294
rect 426986 32378 427222 32614
rect 427306 32378 427542 32614
rect 426986 32058 427222 32294
rect 427306 32058 427542 32294
rect 408986 -6342 409222 -6106
rect 409306 -6342 409542 -6106
rect 408986 -6662 409222 -6426
rect 409306 -6662 409542 -6426
rect 433826 704602 434062 704838
rect 434146 704602 434382 704838
rect 433826 704282 434062 704518
rect 434146 704282 434382 704518
rect 433826 687218 434062 687454
rect 434146 687218 434382 687454
rect 433826 686898 434062 687134
rect 434146 686898 434382 687134
rect 433826 651218 434062 651454
rect 434146 651218 434382 651454
rect 433826 650898 434062 651134
rect 434146 650898 434382 651134
rect 433826 615218 434062 615454
rect 434146 615218 434382 615454
rect 433826 614898 434062 615134
rect 434146 614898 434382 615134
rect 433826 579218 434062 579454
rect 434146 579218 434382 579454
rect 433826 578898 434062 579134
rect 434146 578898 434382 579134
rect 433826 543218 434062 543454
rect 434146 543218 434382 543454
rect 433826 542898 434062 543134
rect 434146 542898 434382 543134
rect 433826 507218 434062 507454
rect 434146 507218 434382 507454
rect 433826 506898 434062 507134
rect 434146 506898 434382 507134
rect 433826 471218 434062 471454
rect 434146 471218 434382 471454
rect 433826 470898 434062 471134
rect 434146 470898 434382 471134
rect 433826 435218 434062 435454
rect 434146 435218 434382 435454
rect 433826 434898 434062 435134
rect 434146 434898 434382 435134
rect 433826 399218 434062 399454
rect 434146 399218 434382 399454
rect 433826 398898 434062 399134
rect 434146 398898 434382 399134
rect 433826 363218 434062 363454
rect 434146 363218 434382 363454
rect 433826 362898 434062 363134
rect 434146 362898 434382 363134
rect 433826 327218 434062 327454
rect 434146 327218 434382 327454
rect 433826 326898 434062 327134
rect 434146 326898 434382 327134
rect 433826 291218 434062 291454
rect 434146 291218 434382 291454
rect 433826 290898 434062 291134
rect 434146 290898 434382 291134
rect 433826 255218 434062 255454
rect 434146 255218 434382 255454
rect 433826 254898 434062 255134
rect 434146 254898 434382 255134
rect 433826 219218 434062 219454
rect 434146 219218 434382 219454
rect 433826 218898 434062 219134
rect 434146 218898 434382 219134
rect 433826 183218 434062 183454
rect 434146 183218 434382 183454
rect 433826 182898 434062 183134
rect 434146 182898 434382 183134
rect 433826 147218 434062 147454
rect 434146 147218 434382 147454
rect 433826 146898 434062 147134
rect 434146 146898 434382 147134
rect 433826 111218 434062 111454
rect 434146 111218 434382 111454
rect 433826 110898 434062 111134
rect 434146 110898 434382 111134
rect 433826 75218 434062 75454
rect 434146 75218 434382 75454
rect 433826 74898 434062 75134
rect 434146 74898 434382 75134
rect 433826 39218 434062 39454
rect 434146 39218 434382 39454
rect 433826 38898 434062 39134
rect 434146 38898 434382 39134
rect 433826 3218 434062 3454
rect 434146 3218 434382 3454
rect 433826 2898 434062 3134
rect 434146 2898 434382 3134
rect 433826 -582 434062 -346
rect 434146 -582 434382 -346
rect 433826 -902 434062 -666
rect 434146 -902 434382 -666
rect 437546 690938 437782 691174
rect 437866 690938 438102 691174
rect 437546 690618 437782 690854
rect 437866 690618 438102 690854
rect 437546 654938 437782 655174
rect 437866 654938 438102 655174
rect 437546 654618 437782 654854
rect 437866 654618 438102 654854
rect 437546 618938 437782 619174
rect 437866 618938 438102 619174
rect 437546 618618 437782 618854
rect 437866 618618 438102 618854
rect 437546 582938 437782 583174
rect 437866 582938 438102 583174
rect 437546 582618 437782 582854
rect 437866 582618 438102 582854
rect 437546 546938 437782 547174
rect 437866 546938 438102 547174
rect 437546 546618 437782 546854
rect 437866 546618 438102 546854
rect 437546 510938 437782 511174
rect 437866 510938 438102 511174
rect 437546 510618 437782 510854
rect 437866 510618 438102 510854
rect 437546 474938 437782 475174
rect 437866 474938 438102 475174
rect 437546 474618 437782 474854
rect 437866 474618 438102 474854
rect 437546 438938 437782 439174
rect 437866 438938 438102 439174
rect 437546 438618 437782 438854
rect 437866 438618 438102 438854
rect 437546 402938 437782 403174
rect 437866 402938 438102 403174
rect 437546 402618 437782 402854
rect 437866 402618 438102 402854
rect 437546 366938 437782 367174
rect 437866 366938 438102 367174
rect 437546 366618 437782 366854
rect 437866 366618 438102 366854
rect 437546 330938 437782 331174
rect 437866 330938 438102 331174
rect 437546 330618 437782 330854
rect 437866 330618 438102 330854
rect 437546 294938 437782 295174
rect 437866 294938 438102 295174
rect 437546 294618 437782 294854
rect 437866 294618 438102 294854
rect 437546 258938 437782 259174
rect 437866 258938 438102 259174
rect 437546 258618 437782 258854
rect 437866 258618 438102 258854
rect 437546 222938 437782 223174
rect 437866 222938 438102 223174
rect 437546 222618 437782 222854
rect 437866 222618 438102 222854
rect 437546 186938 437782 187174
rect 437866 186938 438102 187174
rect 437546 186618 437782 186854
rect 437866 186618 438102 186854
rect 437546 150938 437782 151174
rect 437866 150938 438102 151174
rect 437546 150618 437782 150854
rect 437866 150618 438102 150854
rect 437546 114938 437782 115174
rect 437866 114938 438102 115174
rect 437546 114618 437782 114854
rect 437866 114618 438102 114854
rect 437546 78938 437782 79174
rect 437866 78938 438102 79174
rect 437546 78618 437782 78854
rect 437866 78618 438102 78854
rect 437546 42938 437782 43174
rect 437866 42938 438102 43174
rect 437546 42618 437782 42854
rect 437866 42618 438102 42854
rect 437546 6938 437782 7174
rect 437866 6938 438102 7174
rect 437546 6618 437782 6854
rect 437866 6618 438102 6854
rect 437546 -2502 437782 -2266
rect 437866 -2502 438102 -2266
rect 437546 -2822 437782 -2586
rect 437866 -2822 438102 -2586
rect 441266 694658 441502 694894
rect 441586 694658 441822 694894
rect 441266 694338 441502 694574
rect 441586 694338 441822 694574
rect 441266 658658 441502 658894
rect 441586 658658 441822 658894
rect 441266 658338 441502 658574
rect 441586 658338 441822 658574
rect 441266 622658 441502 622894
rect 441586 622658 441822 622894
rect 441266 622338 441502 622574
rect 441586 622338 441822 622574
rect 441266 586658 441502 586894
rect 441586 586658 441822 586894
rect 441266 586338 441502 586574
rect 441586 586338 441822 586574
rect 441266 550658 441502 550894
rect 441586 550658 441822 550894
rect 441266 550338 441502 550574
rect 441586 550338 441822 550574
rect 441266 514658 441502 514894
rect 441586 514658 441822 514894
rect 441266 514338 441502 514574
rect 441586 514338 441822 514574
rect 441266 478658 441502 478894
rect 441586 478658 441822 478894
rect 441266 478338 441502 478574
rect 441586 478338 441822 478574
rect 441266 442658 441502 442894
rect 441586 442658 441822 442894
rect 441266 442338 441502 442574
rect 441586 442338 441822 442574
rect 441266 406658 441502 406894
rect 441586 406658 441822 406894
rect 441266 406338 441502 406574
rect 441586 406338 441822 406574
rect 441266 370658 441502 370894
rect 441586 370658 441822 370894
rect 441266 370338 441502 370574
rect 441586 370338 441822 370574
rect 441266 334658 441502 334894
rect 441586 334658 441822 334894
rect 441266 334338 441502 334574
rect 441586 334338 441822 334574
rect 441266 298658 441502 298894
rect 441586 298658 441822 298894
rect 441266 298338 441502 298574
rect 441586 298338 441822 298574
rect 441266 262658 441502 262894
rect 441586 262658 441822 262894
rect 441266 262338 441502 262574
rect 441586 262338 441822 262574
rect 441266 226658 441502 226894
rect 441586 226658 441822 226894
rect 441266 226338 441502 226574
rect 441586 226338 441822 226574
rect 441266 190658 441502 190894
rect 441586 190658 441822 190894
rect 441266 190338 441502 190574
rect 441586 190338 441822 190574
rect 441266 154658 441502 154894
rect 441586 154658 441822 154894
rect 441266 154338 441502 154574
rect 441586 154338 441822 154574
rect 441266 118658 441502 118894
rect 441586 118658 441822 118894
rect 441266 118338 441502 118574
rect 441586 118338 441822 118574
rect 441266 82658 441502 82894
rect 441586 82658 441822 82894
rect 441266 82338 441502 82574
rect 441586 82338 441822 82574
rect 441266 46658 441502 46894
rect 441586 46658 441822 46894
rect 441266 46338 441502 46574
rect 441586 46338 441822 46574
rect 441266 10658 441502 10894
rect 441586 10658 441822 10894
rect 441266 10338 441502 10574
rect 441586 10338 441822 10574
rect 441266 -4422 441502 -4186
rect 441586 -4422 441822 -4186
rect 441266 -4742 441502 -4506
rect 441586 -4742 441822 -4506
rect 462986 711322 463222 711558
rect 463306 711322 463542 711558
rect 462986 711002 463222 711238
rect 463306 711002 463542 711238
rect 459266 709402 459502 709638
rect 459586 709402 459822 709638
rect 459266 709082 459502 709318
rect 459586 709082 459822 709318
rect 455546 707482 455782 707718
rect 455866 707482 456102 707718
rect 455546 707162 455782 707398
rect 455866 707162 456102 707398
rect 444986 698378 445222 698614
rect 445306 698378 445542 698614
rect 444986 698058 445222 698294
rect 445306 698058 445542 698294
rect 444986 662378 445222 662614
rect 445306 662378 445542 662614
rect 444986 662058 445222 662294
rect 445306 662058 445542 662294
rect 444986 626378 445222 626614
rect 445306 626378 445542 626614
rect 444986 626058 445222 626294
rect 445306 626058 445542 626294
rect 444986 590378 445222 590614
rect 445306 590378 445542 590614
rect 444986 590058 445222 590294
rect 445306 590058 445542 590294
rect 444986 554378 445222 554614
rect 445306 554378 445542 554614
rect 444986 554058 445222 554294
rect 445306 554058 445542 554294
rect 444986 518378 445222 518614
rect 445306 518378 445542 518614
rect 444986 518058 445222 518294
rect 445306 518058 445542 518294
rect 444986 482378 445222 482614
rect 445306 482378 445542 482614
rect 444986 482058 445222 482294
rect 445306 482058 445542 482294
rect 444986 446378 445222 446614
rect 445306 446378 445542 446614
rect 444986 446058 445222 446294
rect 445306 446058 445542 446294
rect 444986 410378 445222 410614
rect 445306 410378 445542 410614
rect 444986 410058 445222 410294
rect 445306 410058 445542 410294
rect 444986 374378 445222 374614
rect 445306 374378 445542 374614
rect 444986 374058 445222 374294
rect 445306 374058 445542 374294
rect 444986 338378 445222 338614
rect 445306 338378 445542 338614
rect 444986 338058 445222 338294
rect 445306 338058 445542 338294
rect 444986 302378 445222 302614
rect 445306 302378 445542 302614
rect 444986 302058 445222 302294
rect 445306 302058 445542 302294
rect 444986 266378 445222 266614
rect 445306 266378 445542 266614
rect 444986 266058 445222 266294
rect 445306 266058 445542 266294
rect 444986 230378 445222 230614
rect 445306 230378 445542 230614
rect 444986 230058 445222 230294
rect 445306 230058 445542 230294
rect 444986 194378 445222 194614
rect 445306 194378 445542 194614
rect 444986 194058 445222 194294
rect 445306 194058 445542 194294
rect 444986 158378 445222 158614
rect 445306 158378 445542 158614
rect 444986 158058 445222 158294
rect 445306 158058 445542 158294
rect 444986 122378 445222 122614
rect 445306 122378 445542 122614
rect 444986 122058 445222 122294
rect 445306 122058 445542 122294
rect 444986 86378 445222 86614
rect 445306 86378 445542 86614
rect 444986 86058 445222 86294
rect 445306 86058 445542 86294
rect 444986 50378 445222 50614
rect 445306 50378 445542 50614
rect 444986 50058 445222 50294
rect 445306 50058 445542 50294
rect 444986 14378 445222 14614
rect 445306 14378 445542 14614
rect 444986 14058 445222 14294
rect 445306 14058 445542 14294
rect 426986 -7302 427222 -7066
rect 427306 -7302 427542 -7066
rect 426986 -7622 427222 -7386
rect 427306 -7622 427542 -7386
rect 451826 705562 452062 705798
rect 452146 705562 452382 705798
rect 451826 705242 452062 705478
rect 452146 705242 452382 705478
rect 451826 669218 452062 669454
rect 452146 669218 452382 669454
rect 451826 668898 452062 669134
rect 452146 668898 452382 669134
rect 451826 633218 452062 633454
rect 452146 633218 452382 633454
rect 451826 632898 452062 633134
rect 452146 632898 452382 633134
rect 451826 597218 452062 597454
rect 452146 597218 452382 597454
rect 451826 596898 452062 597134
rect 452146 596898 452382 597134
rect 451826 561218 452062 561454
rect 452146 561218 452382 561454
rect 451826 560898 452062 561134
rect 452146 560898 452382 561134
rect 451826 525218 452062 525454
rect 452146 525218 452382 525454
rect 451826 524898 452062 525134
rect 452146 524898 452382 525134
rect 451826 489218 452062 489454
rect 452146 489218 452382 489454
rect 451826 488898 452062 489134
rect 452146 488898 452382 489134
rect 451826 453218 452062 453454
rect 452146 453218 452382 453454
rect 451826 452898 452062 453134
rect 452146 452898 452382 453134
rect 451826 417218 452062 417454
rect 452146 417218 452382 417454
rect 451826 416898 452062 417134
rect 452146 416898 452382 417134
rect 451826 381218 452062 381454
rect 452146 381218 452382 381454
rect 451826 380898 452062 381134
rect 452146 380898 452382 381134
rect 451826 345218 452062 345454
rect 452146 345218 452382 345454
rect 451826 344898 452062 345134
rect 452146 344898 452382 345134
rect 451826 309218 452062 309454
rect 452146 309218 452382 309454
rect 451826 308898 452062 309134
rect 452146 308898 452382 309134
rect 451826 273218 452062 273454
rect 452146 273218 452382 273454
rect 451826 272898 452062 273134
rect 452146 272898 452382 273134
rect 451826 237218 452062 237454
rect 452146 237218 452382 237454
rect 451826 236898 452062 237134
rect 452146 236898 452382 237134
rect 451826 201218 452062 201454
rect 452146 201218 452382 201454
rect 451826 200898 452062 201134
rect 452146 200898 452382 201134
rect 451826 165218 452062 165454
rect 452146 165218 452382 165454
rect 451826 164898 452062 165134
rect 452146 164898 452382 165134
rect 451826 129218 452062 129454
rect 452146 129218 452382 129454
rect 451826 128898 452062 129134
rect 452146 128898 452382 129134
rect 451826 93218 452062 93454
rect 452146 93218 452382 93454
rect 451826 92898 452062 93134
rect 452146 92898 452382 93134
rect 451826 57218 452062 57454
rect 452146 57218 452382 57454
rect 451826 56898 452062 57134
rect 452146 56898 452382 57134
rect 451826 21218 452062 21454
rect 452146 21218 452382 21454
rect 451826 20898 452062 21134
rect 452146 20898 452382 21134
rect 451826 -1542 452062 -1306
rect 452146 -1542 452382 -1306
rect 451826 -1862 452062 -1626
rect 452146 -1862 452382 -1626
rect 455546 672938 455782 673174
rect 455866 672938 456102 673174
rect 455546 672618 455782 672854
rect 455866 672618 456102 672854
rect 455546 636938 455782 637174
rect 455866 636938 456102 637174
rect 455546 636618 455782 636854
rect 455866 636618 456102 636854
rect 455546 600938 455782 601174
rect 455866 600938 456102 601174
rect 455546 600618 455782 600854
rect 455866 600618 456102 600854
rect 455546 564938 455782 565174
rect 455866 564938 456102 565174
rect 455546 564618 455782 564854
rect 455866 564618 456102 564854
rect 455546 528938 455782 529174
rect 455866 528938 456102 529174
rect 455546 528618 455782 528854
rect 455866 528618 456102 528854
rect 455546 492938 455782 493174
rect 455866 492938 456102 493174
rect 455546 492618 455782 492854
rect 455866 492618 456102 492854
rect 455546 456938 455782 457174
rect 455866 456938 456102 457174
rect 455546 456618 455782 456854
rect 455866 456618 456102 456854
rect 455546 420938 455782 421174
rect 455866 420938 456102 421174
rect 455546 420618 455782 420854
rect 455866 420618 456102 420854
rect 455546 384938 455782 385174
rect 455866 384938 456102 385174
rect 455546 384618 455782 384854
rect 455866 384618 456102 384854
rect 455546 348938 455782 349174
rect 455866 348938 456102 349174
rect 455546 348618 455782 348854
rect 455866 348618 456102 348854
rect 455546 312938 455782 313174
rect 455866 312938 456102 313174
rect 455546 312618 455782 312854
rect 455866 312618 456102 312854
rect 455546 276938 455782 277174
rect 455866 276938 456102 277174
rect 455546 276618 455782 276854
rect 455866 276618 456102 276854
rect 455546 240938 455782 241174
rect 455866 240938 456102 241174
rect 455546 240618 455782 240854
rect 455866 240618 456102 240854
rect 455546 204938 455782 205174
rect 455866 204938 456102 205174
rect 455546 204618 455782 204854
rect 455866 204618 456102 204854
rect 455546 168938 455782 169174
rect 455866 168938 456102 169174
rect 455546 168618 455782 168854
rect 455866 168618 456102 168854
rect 455546 132938 455782 133174
rect 455866 132938 456102 133174
rect 455546 132618 455782 132854
rect 455866 132618 456102 132854
rect 455546 96938 455782 97174
rect 455866 96938 456102 97174
rect 455546 96618 455782 96854
rect 455866 96618 456102 96854
rect 455546 60938 455782 61174
rect 455866 60938 456102 61174
rect 455546 60618 455782 60854
rect 455866 60618 456102 60854
rect 455546 24938 455782 25174
rect 455866 24938 456102 25174
rect 455546 24618 455782 24854
rect 455866 24618 456102 24854
rect 455546 -3462 455782 -3226
rect 455866 -3462 456102 -3226
rect 455546 -3782 455782 -3546
rect 455866 -3782 456102 -3546
rect 459266 676658 459502 676894
rect 459586 676658 459822 676894
rect 459266 676338 459502 676574
rect 459586 676338 459822 676574
rect 459266 640658 459502 640894
rect 459586 640658 459822 640894
rect 459266 640338 459502 640574
rect 459586 640338 459822 640574
rect 459266 604658 459502 604894
rect 459586 604658 459822 604894
rect 459266 604338 459502 604574
rect 459586 604338 459822 604574
rect 459266 568658 459502 568894
rect 459586 568658 459822 568894
rect 459266 568338 459502 568574
rect 459586 568338 459822 568574
rect 459266 532658 459502 532894
rect 459586 532658 459822 532894
rect 459266 532338 459502 532574
rect 459586 532338 459822 532574
rect 459266 496658 459502 496894
rect 459586 496658 459822 496894
rect 459266 496338 459502 496574
rect 459586 496338 459822 496574
rect 459266 460658 459502 460894
rect 459586 460658 459822 460894
rect 459266 460338 459502 460574
rect 459586 460338 459822 460574
rect 459266 424658 459502 424894
rect 459586 424658 459822 424894
rect 459266 424338 459502 424574
rect 459586 424338 459822 424574
rect 459266 388658 459502 388894
rect 459586 388658 459822 388894
rect 459266 388338 459502 388574
rect 459586 388338 459822 388574
rect 459266 352658 459502 352894
rect 459586 352658 459822 352894
rect 459266 352338 459502 352574
rect 459586 352338 459822 352574
rect 459266 316658 459502 316894
rect 459586 316658 459822 316894
rect 459266 316338 459502 316574
rect 459586 316338 459822 316574
rect 459266 280658 459502 280894
rect 459586 280658 459822 280894
rect 459266 280338 459502 280574
rect 459586 280338 459822 280574
rect 459266 244658 459502 244894
rect 459586 244658 459822 244894
rect 459266 244338 459502 244574
rect 459586 244338 459822 244574
rect 459266 208658 459502 208894
rect 459586 208658 459822 208894
rect 459266 208338 459502 208574
rect 459586 208338 459822 208574
rect 459266 172658 459502 172894
rect 459586 172658 459822 172894
rect 459266 172338 459502 172574
rect 459586 172338 459822 172574
rect 459266 136658 459502 136894
rect 459586 136658 459822 136894
rect 459266 136338 459502 136574
rect 459586 136338 459822 136574
rect 459266 100658 459502 100894
rect 459586 100658 459822 100894
rect 459266 100338 459502 100574
rect 459586 100338 459822 100574
rect 459266 64658 459502 64894
rect 459586 64658 459822 64894
rect 459266 64338 459502 64574
rect 459586 64338 459822 64574
rect 459266 28658 459502 28894
rect 459586 28658 459822 28894
rect 459266 28338 459502 28574
rect 459586 28338 459822 28574
rect 459266 -5382 459502 -5146
rect 459586 -5382 459822 -5146
rect 459266 -5702 459502 -5466
rect 459586 -5702 459822 -5466
rect 480986 710362 481222 710598
rect 481306 710362 481542 710598
rect 480986 710042 481222 710278
rect 481306 710042 481542 710278
rect 477266 708442 477502 708678
rect 477586 708442 477822 708678
rect 477266 708122 477502 708358
rect 477586 708122 477822 708358
rect 473546 706522 473782 706758
rect 473866 706522 474102 706758
rect 473546 706202 473782 706438
rect 473866 706202 474102 706438
rect 462986 680378 463222 680614
rect 463306 680378 463542 680614
rect 462986 680058 463222 680294
rect 463306 680058 463542 680294
rect 462986 644378 463222 644614
rect 463306 644378 463542 644614
rect 462986 644058 463222 644294
rect 463306 644058 463542 644294
rect 462986 608378 463222 608614
rect 463306 608378 463542 608614
rect 462986 608058 463222 608294
rect 463306 608058 463542 608294
rect 462986 572378 463222 572614
rect 463306 572378 463542 572614
rect 462986 572058 463222 572294
rect 463306 572058 463542 572294
rect 462986 536378 463222 536614
rect 463306 536378 463542 536614
rect 462986 536058 463222 536294
rect 463306 536058 463542 536294
rect 462986 500378 463222 500614
rect 463306 500378 463542 500614
rect 462986 500058 463222 500294
rect 463306 500058 463542 500294
rect 462986 464378 463222 464614
rect 463306 464378 463542 464614
rect 462986 464058 463222 464294
rect 463306 464058 463542 464294
rect 462986 428378 463222 428614
rect 463306 428378 463542 428614
rect 462986 428058 463222 428294
rect 463306 428058 463542 428294
rect 462986 392378 463222 392614
rect 463306 392378 463542 392614
rect 462986 392058 463222 392294
rect 463306 392058 463542 392294
rect 462986 356378 463222 356614
rect 463306 356378 463542 356614
rect 462986 356058 463222 356294
rect 463306 356058 463542 356294
rect 462986 320378 463222 320614
rect 463306 320378 463542 320614
rect 462986 320058 463222 320294
rect 463306 320058 463542 320294
rect 462986 284378 463222 284614
rect 463306 284378 463542 284614
rect 462986 284058 463222 284294
rect 463306 284058 463542 284294
rect 462986 248378 463222 248614
rect 463306 248378 463542 248614
rect 462986 248058 463222 248294
rect 463306 248058 463542 248294
rect 462986 212378 463222 212614
rect 463306 212378 463542 212614
rect 462986 212058 463222 212294
rect 463306 212058 463542 212294
rect 462986 176378 463222 176614
rect 463306 176378 463542 176614
rect 462986 176058 463222 176294
rect 463306 176058 463542 176294
rect 462986 140378 463222 140614
rect 463306 140378 463542 140614
rect 462986 140058 463222 140294
rect 463306 140058 463542 140294
rect 462986 104378 463222 104614
rect 463306 104378 463542 104614
rect 462986 104058 463222 104294
rect 463306 104058 463542 104294
rect 462986 68378 463222 68614
rect 463306 68378 463542 68614
rect 462986 68058 463222 68294
rect 463306 68058 463542 68294
rect 462986 32378 463222 32614
rect 463306 32378 463542 32614
rect 462986 32058 463222 32294
rect 463306 32058 463542 32294
rect 444986 -6342 445222 -6106
rect 445306 -6342 445542 -6106
rect 444986 -6662 445222 -6426
rect 445306 -6662 445542 -6426
rect 469826 704602 470062 704838
rect 470146 704602 470382 704838
rect 469826 704282 470062 704518
rect 470146 704282 470382 704518
rect 469826 687218 470062 687454
rect 470146 687218 470382 687454
rect 469826 686898 470062 687134
rect 470146 686898 470382 687134
rect 469826 651218 470062 651454
rect 470146 651218 470382 651454
rect 469826 650898 470062 651134
rect 470146 650898 470382 651134
rect 469826 615218 470062 615454
rect 470146 615218 470382 615454
rect 469826 614898 470062 615134
rect 470146 614898 470382 615134
rect 469826 579218 470062 579454
rect 470146 579218 470382 579454
rect 469826 578898 470062 579134
rect 470146 578898 470382 579134
rect 469826 543218 470062 543454
rect 470146 543218 470382 543454
rect 469826 542898 470062 543134
rect 470146 542898 470382 543134
rect 469826 507218 470062 507454
rect 470146 507218 470382 507454
rect 469826 506898 470062 507134
rect 470146 506898 470382 507134
rect 469826 471218 470062 471454
rect 470146 471218 470382 471454
rect 469826 470898 470062 471134
rect 470146 470898 470382 471134
rect 469826 435218 470062 435454
rect 470146 435218 470382 435454
rect 469826 434898 470062 435134
rect 470146 434898 470382 435134
rect 469826 399218 470062 399454
rect 470146 399218 470382 399454
rect 469826 398898 470062 399134
rect 470146 398898 470382 399134
rect 469826 363218 470062 363454
rect 470146 363218 470382 363454
rect 469826 362898 470062 363134
rect 470146 362898 470382 363134
rect 469826 327218 470062 327454
rect 470146 327218 470382 327454
rect 469826 326898 470062 327134
rect 470146 326898 470382 327134
rect 469826 291218 470062 291454
rect 470146 291218 470382 291454
rect 469826 290898 470062 291134
rect 470146 290898 470382 291134
rect 469826 255218 470062 255454
rect 470146 255218 470382 255454
rect 469826 254898 470062 255134
rect 470146 254898 470382 255134
rect 469826 219218 470062 219454
rect 470146 219218 470382 219454
rect 469826 218898 470062 219134
rect 470146 218898 470382 219134
rect 469826 183218 470062 183454
rect 470146 183218 470382 183454
rect 469826 182898 470062 183134
rect 470146 182898 470382 183134
rect 469826 147218 470062 147454
rect 470146 147218 470382 147454
rect 469826 146898 470062 147134
rect 470146 146898 470382 147134
rect 469826 111218 470062 111454
rect 470146 111218 470382 111454
rect 469826 110898 470062 111134
rect 470146 110898 470382 111134
rect 469826 75218 470062 75454
rect 470146 75218 470382 75454
rect 469826 74898 470062 75134
rect 470146 74898 470382 75134
rect 469826 39218 470062 39454
rect 470146 39218 470382 39454
rect 469826 38898 470062 39134
rect 470146 38898 470382 39134
rect 469826 3218 470062 3454
rect 470146 3218 470382 3454
rect 469826 2898 470062 3134
rect 470146 2898 470382 3134
rect 469826 -582 470062 -346
rect 470146 -582 470382 -346
rect 469826 -902 470062 -666
rect 470146 -902 470382 -666
rect 473546 690938 473782 691174
rect 473866 690938 474102 691174
rect 473546 690618 473782 690854
rect 473866 690618 474102 690854
rect 473546 654938 473782 655174
rect 473866 654938 474102 655174
rect 473546 654618 473782 654854
rect 473866 654618 474102 654854
rect 473546 618938 473782 619174
rect 473866 618938 474102 619174
rect 473546 618618 473782 618854
rect 473866 618618 474102 618854
rect 473546 582938 473782 583174
rect 473866 582938 474102 583174
rect 473546 582618 473782 582854
rect 473866 582618 474102 582854
rect 473546 546938 473782 547174
rect 473866 546938 474102 547174
rect 473546 546618 473782 546854
rect 473866 546618 474102 546854
rect 473546 510938 473782 511174
rect 473866 510938 474102 511174
rect 473546 510618 473782 510854
rect 473866 510618 474102 510854
rect 473546 474938 473782 475174
rect 473866 474938 474102 475174
rect 473546 474618 473782 474854
rect 473866 474618 474102 474854
rect 473546 438938 473782 439174
rect 473866 438938 474102 439174
rect 473546 438618 473782 438854
rect 473866 438618 474102 438854
rect 473546 402938 473782 403174
rect 473866 402938 474102 403174
rect 473546 402618 473782 402854
rect 473866 402618 474102 402854
rect 473546 366938 473782 367174
rect 473866 366938 474102 367174
rect 473546 366618 473782 366854
rect 473866 366618 474102 366854
rect 473546 330938 473782 331174
rect 473866 330938 474102 331174
rect 473546 330618 473782 330854
rect 473866 330618 474102 330854
rect 473546 294938 473782 295174
rect 473866 294938 474102 295174
rect 473546 294618 473782 294854
rect 473866 294618 474102 294854
rect 473546 258938 473782 259174
rect 473866 258938 474102 259174
rect 473546 258618 473782 258854
rect 473866 258618 474102 258854
rect 473546 222938 473782 223174
rect 473866 222938 474102 223174
rect 473546 222618 473782 222854
rect 473866 222618 474102 222854
rect 473546 186938 473782 187174
rect 473866 186938 474102 187174
rect 473546 186618 473782 186854
rect 473866 186618 474102 186854
rect 473546 150938 473782 151174
rect 473866 150938 474102 151174
rect 473546 150618 473782 150854
rect 473866 150618 474102 150854
rect 473546 114938 473782 115174
rect 473866 114938 474102 115174
rect 473546 114618 473782 114854
rect 473866 114618 474102 114854
rect 473546 78938 473782 79174
rect 473866 78938 474102 79174
rect 473546 78618 473782 78854
rect 473866 78618 474102 78854
rect 473546 42938 473782 43174
rect 473866 42938 474102 43174
rect 473546 42618 473782 42854
rect 473866 42618 474102 42854
rect 473546 6938 473782 7174
rect 473866 6938 474102 7174
rect 473546 6618 473782 6854
rect 473866 6618 474102 6854
rect 473546 -2502 473782 -2266
rect 473866 -2502 474102 -2266
rect 473546 -2822 473782 -2586
rect 473866 -2822 474102 -2586
rect 477266 694658 477502 694894
rect 477586 694658 477822 694894
rect 477266 694338 477502 694574
rect 477586 694338 477822 694574
rect 477266 658658 477502 658894
rect 477586 658658 477822 658894
rect 477266 658338 477502 658574
rect 477586 658338 477822 658574
rect 477266 622658 477502 622894
rect 477586 622658 477822 622894
rect 477266 622338 477502 622574
rect 477586 622338 477822 622574
rect 477266 586658 477502 586894
rect 477586 586658 477822 586894
rect 477266 586338 477502 586574
rect 477586 586338 477822 586574
rect 477266 550658 477502 550894
rect 477586 550658 477822 550894
rect 477266 550338 477502 550574
rect 477586 550338 477822 550574
rect 477266 514658 477502 514894
rect 477586 514658 477822 514894
rect 477266 514338 477502 514574
rect 477586 514338 477822 514574
rect 477266 478658 477502 478894
rect 477586 478658 477822 478894
rect 477266 478338 477502 478574
rect 477586 478338 477822 478574
rect 477266 442658 477502 442894
rect 477586 442658 477822 442894
rect 477266 442338 477502 442574
rect 477586 442338 477822 442574
rect 477266 406658 477502 406894
rect 477586 406658 477822 406894
rect 477266 406338 477502 406574
rect 477586 406338 477822 406574
rect 477266 370658 477502 370894
rect 477586 370658 477822 370894
rect 477266 370338 477502 370574
rect 477586 370338 477822 370574
rect 477266 334658 477502 334894
rect 477586 334658 477822 334894
rect 477266 334338 477502 334574
rect 477586 334338 477822 334574
rect 477266 298658 477502 298894
rect 477586 298658 477822 298894
rect 477266 298338 477502 298574
rect 477586 298338 477822 298574
rect 477266 262658 477502 262894
rect 477586 262658 477822 262894
rect 477266 262338 477502 262574
rect 477586 262338 477822 262574
rect 477266 226658 477502 226894
rect 477586 226658 477822 226894
rect 477266 226338 477502 226574
rect 477586 226338 477822 226574
rect 477266 190658 477502 190894
rect 477586 190658 477822 190894
rect 477266 190338 477502 190574
rect 477586 190338 477822 190574
rect 477266 154658 477502 154894
rect 477586 154658 477822 154894
rect 477266 154338 477502 154574
rect 477586 154338 477822 154574
rect 477266 118658 477502 118894
rect 477586 118658 477822 118894
rect 477266 118338 477502 118574
rect 477586 118338 477822 118574
rect 477266 82658 477502 82894
rect 477586 82658 477822 82894
rect 477266 82338 477502 82574
rect 477586 82338 477822 82574
rect 477266 46658 477502 46894
rect 477586 46658 477822 46894
rect 477266 46338 477502 46574
rect 477586 46338 477822 46574
rect 477266 10658 477502 10894
rect 477586 10658 477822 10894
rect 477266 10338 477502 10574
rect 477586 10338 477822 10574
rect 477266 -4422 477502 -4186
rect 477586 -4422 477822 -4186
rect 477266 -4742 477502 -4506
rect 477586 -4742 477822 -4506
rect 498986 711322 499222 711558
rect 499306 711322 499542 711558
rect 498986 711002 499222 711238
rect 499306 711002 499542 711238
rect 495266 709402 495502 709638
rect 495586 709402 495822 709638
rect 495266 709082 495502 709318
rect 495586 709082 495822 709318
rect 491546 707482 491782 707718
rect 491866 707482 492102 707718
rect 491546 707162 491782 707398
rect 491866 707162 492102 707398
rect 480986 698378 481222 698614
rect 481306 698378 481542 698614
rect 480986 698058 481222 698294
rect 481306 698058 481542 698294
rect 480986 662378 481222 662614
rect 481306 662378 481542 662614
rect 480986 662058 481222 662294
rect 481306 662058 481542 662294
rect 480986 626378 481222 626614
rect 481306 626378 481542 626614
rect 480986 626058 481222 626294
rect 481306 626058 481542 626294
rect 480986 590378 481222 590614
rect 481306 590378 481542 590614
rect 480986 590058 481222 590294
rect 481306 590058 481542 590294
rect 480986 554378 481222 554614
rect 481306 554378 481542 554614
rect 480986 554058 481222 554294
rect 481306 554058 481542 554294
rect 480986 518378 481222 518614
rect 481306 518378 481542 518614
rect 480986 518058 481222 518294
rect 481306 518058 481542 518294
rect 480986 482378 481222 482614
rect 481306 482378 481542 482614
rect 480986 482058 481222 482294
rect 481306 482058 481542 482294
rect 480986 446378 481222 446614
rect 481306 446378 481542 446614
rect 480986 446058 481222 446294
rect 481306 446058 481542 446294
rect 480986 410378 481222 410614
rect 481306 410378 481542 410614
rect 480986 410058 481222 410294
rect 481306 410058 481542 410294
rect 480986 374378 481222 374614
rect 481306 374378 481542 374614
rect 480986 374058 481222 374294
rect 481306 374058 481542 374294
rect 480986 338378 481222 338614
rect 481306 338378 481542 338614
rect 480986 338058 481222 338294
rect 481306 338058 481542 338294
rect 480986 302378 481222 302614
rect 481306 302378 481542 302614
rect 480986 302058 481222 302294
rect 481306 302058 481542 302294
rect 480986 266378 481222 266614
rect 481306 266378 481542 266614
rect 480986 266058 481222 266294
rect 481306 266058 481542 266294
rect 480986 230378 481222 230614
rect 481306 230378 481542 230614
rect 480986 230058 481222 230294
rect 481306 230058 481542 230294
rect 480986 194378 481222 194614
rect 481306 194378 481542 194614
rect 480986 194058 481222 194294
rect 481306 194058 481542 194294
rect 480986 158378 481222 158614
rect 481306 158378 481542 158614
rect 480986 158058 481222 158294
rect 481306 158058 481542 158294
rect 480986 122378 481222 122614
rect 481306 122378 481542 122614
rect 480986 122058 481222 122294
rect 481306 122058 481542 122294
rect 480986 86378 481222 86614
rect 481306 86378 481542 86614
rect 480986 86058 481222 86294
rect 481306 86058 481542 86294
rect 480986 50378 481222 50614
rect 481306 50378 481542 50614
rect 480986 50058 481222 50294
rect 481306 50058 481542 50294
rect 480986 14378 481222 14614
rect 481306 14378 481542 14614
rect 480986 14058 481222 14294
rect 481306 14058 481542 14294
rect 462986 -7302 463222 -7066
rect 463306 -7302 463542 -7066
rect 462986 -7622 463222 -7386
rect 463306 -7622 463542 -7386
rect 487826 705562 488062 705798
rect 488146 705562 488382 705798
rect 487826 705242 488062 705478
rect 488146 705242 488382 705478
rect 487826 669218 488062 669454
rect 488146 669218 488382 669454
rect 487826 668898 488062 669134
rect 488146 668898 488382 669134
rect 487826 633218 488062 633454
rect 488146 633218 488382 633454
rect 487826 632898 488062 633134
rect 488146 632898 488382 633134
rect 487826 597218 488062 597454
rect 488146 597218 488382 597454
rect 487826 596898 488062 597134
rect 488146 596898 488382 597134
rect 487826 561218 488062 561454
rect 488146 561218 488382 561454
rect 487826 560898 488062 561134
rect 488146 560898 488382 561134
rect 487826 525218 488062 525454
rect 488146 525218 488382 525454
rect 487826 524898 488062 525134
rect 488146 524898 488382 525134
rect 487826 489218 488062 489454
rect 488146 489218 488382 489454
rect 487826 488898 488062 489134
rect 488146 488898 488382 489134
rect 487826 453218 488062 453454
rect 488146 453218 488382 453454
rect 487826 452898 488062 453134
rect 488146 452898 488382 453134
rect 487826 417218 488062 417454
rect 488146 417218 488382 417454
rect 487826 416898 488062 417134
rect 488146 416898 488382 417134
rect 487826 381218 488062 381454
rect 488146 381218 488382 381454
rect 487826 380898 488062 381134
rect 488146 380898 488382 381134
rect 487826 345218 488062 345454
rect 488146 345218 488382 345454
rect 487826 344898 488062 345134
rect 488146 344898 488382 345134
rect 487826 309218 488062 309454
rect 488146 309218 488382 309454
rect 487826 308898 488062 309134
rect 488146 308898 488382 309134
rect 487826 273218 488062 273454
rect 488146 273218 488382 273454
rect 487826 272898 488062 273134
rect 488146 272898 488382 273134
rect 487826 237218 488062 237454
rect 488146 237218 488382 237454
rect 487826 236898 488062 237134
rect 488146 236898 488382 237134
rect 487826 201218 488062 201454
rect 488146 201218 488382 201454
rect 487826 200898 488062 201134
rect 488146 200898 488382 201134
rect 487826 165218 488062 165454
rect 488146 165218 488382 165454
rect 487826 164898 488062 165134
rect 488146 164898 488382 165134
rect 487826 129218 488062 129454
rect 488146 129218 488382 129454
rect 487826 128898 488062 129134
rect 488146 128898 488382 129134
rect 487826 93218 488062 93454
rect 488146 93218 488382 93454
rect 487826 92898 488062 93134
rect 488146 92898 488382 93134
rect 487826 57218 488062 57454
rect 488146 57218 488382 57454
rect 487826 56898 488062 57134
rect 488146 56898 488382 57134
rect 487826 21218 488062 21454
rect 488146 21218 488382 21454
rect 487826 20898 488062 21134
rect 488146 20898 488382 21134
rect 487826 -1542 488062 -1306
rect 488146 -1542 488382 -1306
rect 487826 -1862 488062 -1626
rect 488146 -1862 488382 -1626
rect 491546 672938 491782 673174
rect 491866 672938 492102 673174
rect 491546 672618 491782 672854
rect 491866 672618 492102 672854
rect 491546 636938 491782 637174
rect 491866 636938 492102 637174
rect 491546 636618 491782 636854
rect 491866 636618 492102 636854
rect 491546 600938 491782 601174
rect 491866 600938 492102 601174
rect 491546 600618 491782 600854
rect 491866 600618 492102 600854
rect 491546 564938 491782 565174
rect 491866 564938 492102 565174
rect 491546 564618 491782 564854
rect 491866 564618 492102 564854
rect 491546 528938 491782 529174
rect 491866 528938 492102 529174
rect 491546 528618 491782 528854
rect 491866 528618 492102 528854
rect 491546 492938 491782 493174
rect 491866 492938 492102 493174
rect 491546 492618 491782 492854
rect 491866 492618 492102 492854
rect 491546 456938 491782 457174
rect 491866 456938 492102 457174
rect 491546 456618 491782 456854
rect 491866 456618 492102 456854
rect 491546 420938 491782 421174
rect 491866 420938 492102 421174
rect 491546 420618 491782 420854
rect 491866 420618 492102 420854
rect 491546 384938 491782 385174
rect 491866 384938 492102 385174
rect 491546 384618 491782 384854
rect 491866 384618 492102 384854
rect 491546 348938 491782 349174
rect 491866 348938 492102 349174
rect 491546 348618 491782 348854
rect 491866 348618 492102 348854
rect 491546 312938 491782 313174
rect 491866 312938 492102 313174
rect 491546 312618 491782 312854
rect 491866 312618 492102 312854
rect 491546 276938 491782 277174
rect 491866 276938 492102 277174
rect 491546 276618 491782 276854
rect 491866 276618 492102 276854
rect 491546 240938 491782 241174
rect 491866 240938 492102 241174
rect 491546 240618 491782 240854
rect 491866 240618 492102 240854
rect 491546 204938 491782 205174
rect 491866 204938 492102 205174
rect 491546 204618 491782 204854
rect 491866 204618 492102 204854
rect 491546 168938 491782 169174
rect 491866 168938 492102 169174
rect 491546 168618 491782 168854
rect 491866 168618 492102 168854
rect 491546 132938 491782 133174
rect 491866 132938 492102 133174
rect 491546 132618 491782 132854
rect 491866 132618 492102 132854
rect 491546 96938 491782 97174
rect 491866 96938 492102 97174
rect 491546 96618 491782 96854
rect 491866 96618 492102 96854
rect 491546 60938 491782 61174
rect 491866 60938 492102 61174
rect 491546 60618 491782 60854
rect 491866 60618 492102 60854
rect 491546 24938 491782 25174
rect 491866 24938 492102 25174
rect 491546 24618 491782 24854
rect 491866 24618 492102 24854
rect 491546 -3462 491782 -3226
rect 491866 -3462 492102 -3226
rect 491546 -3782 491782 -3546
rect 491866 -3782 492102 -3546
rect 495266 676658 495502 676894
rect 495586 676658 495822 676894
rect 495266 676338 495502 676574
rect 495586 676338 495822 676574
rect 495266 640658 495502 640894
rect 495586 640658 495822 640894
rect 495266 640338 495502 640574
rect 495586 640338 495822 640574
rect 495266 604658 495502 604894
rect 495586 604658 495822 604894
rect 495266 604338 495502 604574
rect 495586 604338 495822 604574
rect 495266 568658 495502 568894
rect 495586 568658 495822 568894
rect 495266 568338 495502 568574
rect 495586 568338 495822 568574
rect 495266 532658 495502 532894
rect 495586 532658 495822 532894
rect 495266 532338 495502 532574
rect 495586 532338 495822 532574
rect 495266 496658 495502 496894
rect 495586 496658 495822 496894
rect 495266 496338 495502 496574
rect 495586 496338 495822 496574
rect 495266 460658 495502 460894
rect 495586 460658 495822 460894
rect 495266 460338 495502 460574
rect 495586 460338 495822 460574
rect 495266 424658 495502 424894
rect 495586 424658 495822 424894
rect 495266 424338 495502 424574
rect 495586 424338 495822 424574
rect 495266 388658 495502 388894
rect 495586 388658 495822 388894
rect 495266 388338 495502 388574
rect 495586 388338 495822 388574
rect 495266 352658 495502 352894
rect 495586 352658 495822 352894
rect 495266 352338 495502 352574
rect 495586 352338 495822 352574
rect 495266 316658 495502 316894
rect 495586 316658 495822 316894
rect 495266 316338 495502 316574
rect 495586 316338 495822 316574
rect 495266 280658 495502 280894
rect 495586 280658 495822 280894
rect 495266 280338 495502 280574
rect 495586 280338 495822 280574
rect 495266 244658 495502 244894
rect 495586 244658 495822 244894
rect 495266 244338 495502 244574
rect 495586 244338 495822 244574
rect 495266 208658 495502 208894
rect 495586 208658 495822 208894
rect 495266 208338 495502 208574
rect 495586 208338 495822 208574
rect 495266 172658 495502 172894
rect 495586 172658 495822 172894
rect 495266 172338 495502 172574
rect 495586 172338 495822 172574
rect 495266 136658 495502 136894
rect 495586 136658 495822 136894
rect 495266 136338 495502 136574
rect 495586 136338 495822 136574
rect 495266 100658 495502 100894
rect 495586 100658 495822 100894
rect 495266 100338 495502 100574
rect 495586 100338 495822 100574
rect 495266 64658 495502 64894
rect 495586 64658 495822 64894
rect 495266 64338 495502 64574
rect 495586 64338 495822 64574
rect 495266 28658 495502 28894
rect 495586 28658 495822 28894
rect 495266 28338 495502 28574
rect 495586 28338 495822 28574
rect 495266 -5382 495502 -5146
rect 495586 -5382 495822 -5146
rect 495266 -5702 495502 -5466
rect 495586 -5702 495822 -5466
rect 516986 710362 517222 710598
rect 517306 710362 517542 710598
rect 516986 710042 517222 710278
rect 517306 710042 517542 710278
rect 513266 708442 513502 708678
rect 513586 708442 513822 708678
rect 513266 708122 513502 708358
rect 513586 708122 513822 708358
rect 509546 706522 509782 706758
rect 509866 706522 510102 706758
rect 509546 706202 509782 706438
rect 509866 706202 510102 706438
rect 498986 680378 499222 680614
rect 499306 680378 499542 680614
rect 498986 680058 499222 680294
rect 499306 680058 499542 680294
rect 498986 644378 499222 644614
rect 499306 644378 499542 644614
rect 498986 644058 499222 644294
rect 499306 644058 499542 644294
rect 498986 608378 499222 608614
rect 499306 608378 499542 608614
rect 498986 608058 499222 608294
rect 499306 608058 499542 608294
rect 498986 572378 499222 572614
rect 499306 572378 499542 572614
rect 498986 572058 499222 572294
rect 499306 572058 499542 572294
rect 498986 536378 499222 536614
rect 499306 536378 499542 536614
rect 498986 536058 499222 536294
rect 499306 536058 499542 536294
rect 498986 500378 499222 500614
rect 499306 500378 499542 500614
rect 498986 500058 499222 500294
rect 499306 500058 499542 500294
rect 498986 464378 499222 464614
rect 499306 464378 499542 464614
rect 498986 464058 499222 464294
rect 499306 464058 499542 464294
rect 498986 428378 499222 428614
rect 499306 428378 499542 428614
rect 498986 428058 499222 428294
rect 499306 428058 499542 428294
rect 498986 392378 499222 392614
rect 499306 392378 499542 392614
rect 498986 392058 499222 392294
rect 499306 392058 499542 392294
rect 498986 356378 499222 356614
rect 499306 356378 499542 356614
rect 498986 356058 499222 356294
rect 499306 356058 499542 356294
rect 498986 320378 499222 320614
rect 499306 320378 499542 320614
rect 498986 320058 499222 320294
rect 499306 320058 499542 320294
rect 498986 284378 499222 284614
rect 499306 284378 499542 284614
rect 498986 284058 499222 284294
rect 499306 284058 499542 284294
rect 498986 248378 499222 248614
rect 499306 248378 499542 248614
rect 498986 248058 499222 248294
rect 499306 248058 499542 248294
rect 498986 212378 499222 212614
rect 499306 212378 499542 212614
rect 498986 212058 499222 212294
rect 499306 212058 499542 212294
rect 498986 176378 499222 176614
rect 499306 176378 499542 176614
rect 498986 176058 499222 176294
rect 499306 176058 499542 176294
rect 498986 140378 499222 140614
rect 499306 140378 499542 140614
rect 498986 140058 499222 140294
rect 499306 140058 499542 140294
rect 498986 104378 499222 104614
rect 499306 104378 499542 104614
rect 498986 104058 499222 104294
rect 499306 104058 499542 104294
rect 498986 68378 499222 68614
rect 499306 68378 499542 68614
rect 498986 68058 499222 68294
rect 499306 68058 499542 68294
rect 498986 32378 499222 32614
rect 499306 32378 499542 32614
rect 498986 32058 499222 32294
rect 499306 32058 499542 32294
rect 480986 -6342 481222 -6106
rect 481306 -6342 481542 -6106
rect 480986 -6662 481222 -6426
rect 481306 -6662 481542 -6426
rect 505826 704602 506062 704838
rect 506146 704602 506382 704838
rect 505826 704282 506062 704518
rect 506146 704282 506382 704518
rect 505826 687218 506062 687454
rect 506146 687218 506382 687454
rect 505826 686898 506062 687134
rect 506146 686898 506382 687134
rect 505826 651218 506062 651454
rect 506146 651218 506382 651454
rect 505826 650898 506062 651134
rect 506146 650898 506382 651134
rect 505826 615218 506062 615454
rect 506146 615218 506382 615454
rect 505826 614898 506062 615134
rect 506146 614898 506382 615134
rect 505826 579218 506062 579454
rect 506146 579218 506382 579454
rect 505826 578898 506062 579134
rect 506146 578898 506382 579134
rect 505826 543218 506062 543454
rect 506146 543218 506382 543454
rect 505826 542898 506062 543134
rect 506146 542898 506382 543134
rect 505826 507218 506062 507454
rect 506146 507218 506382 507454
rect 505826 506898 506062 507134
rect 506146 506898 506382 507134
rect 505826 471218 506062 471454
rect 506146 471218 506382 471454
rect 505826 470898 506062 471134
rect 506146 470898 506382 471134
rect 505826 435218 506062 435454
rect 506146 435218 506382 435454
rect 505826 434898 506062 435134
rect 506146 434898 506382 435134
rect 505826 399218 506062 399454
rect 506146 399218 506382 399454
rect 505826 398898 506062 399134
rect 506146 398898 506382 399134
rect 505826 363218 506062 363454
rect 506146 363218 506382 363454
rect 505826 362898 506062 363134
rect 506146 362898 506382 363134
rect 505826 327218 506062 327454
rect 506146 327218 506382 327454
rect 505826 326898 506062 327134
rect 506146 326898 506382 327134
rect 505826 291218 506062 291454
rect 506146 291218 506382 291454
rect 505826 290898 506062 291134
rect 506146 290898 506382 291134
rect 505826 255218 506062 255454
rect 506146 255218 506382 255454
rect 505826 254898 506062 255134
rect 506146 254898 506382 255134
rect 505826 219218 506062 219454
rect 506146 219218 506382 219454
rect 505826 218898 506062 219134
rect 506146 218898 506382 219134
rect 505826 183218 506062 183454
rect 506146 183218 506382 183454
rect 505826 182898 506062 183134
rect 506146 182898 506382 183134
rect 505826 147218 506062 147454
rect 506146 147218 506382 147454
rect 505826 146898 506062 147134
rect 506146 146898 506382 147134
rect 505826 111218 506062 111454
rect 506146 111218 506382 111454
rect 505826 110898 506062 111134
rect 506146 110898 506382 111134
rect 505826 75218 506062 75454
rect 506146 75218 506382 75454
rect 505826 74898 506062 75134
rect 506146 74898 506382 75134
rect 505826 39218 506062 39454
rect 506146 39218 506382 39454
rect 505826 38898 506062 39134
rect 506146 38898 506382 39134
rect 505826 3218 506062 3454
rect 506146 3218 506382 3454
rect 505826 2898 506062 3134
rect 506146 2898 506382 3134
rect 505826 -582 506062 -346
rect 506146 -582 506382 -346
rect 505826 -902 506062 -666
rect 506146 -902 506382 -666
rect 509546 690938 509782 691174
rect 509866 690938 510102 691174
rect 509546 690618 509782 690854
rect 509866 690618 510102 690854
rect 509546 654938 509782 655174
rect 509866 654938 510102 655174
rect 509546 654618 509782 654854
rect 509866 654618 510102 654854
rect 509546 618938 509782 619174
rect 509866 618938 510102 619174
rect 509546 618618 509782 618854
rect 509866 618618 510102 618854
rect 509546 582938 509782 583174
rect 509866 582938 510102 583174
rect 509546 582618 509782 582854
rect 509866 582618 510102 582854
rect 509546 546938 509782 547174
rect 509866 546938 510102 547174
rect 509546 546618 509782 546854
rect 509866 546618 510102 546854
rect 509546 510938 509782 511174
rect 509866 510938 510102 511174
rect 509546 510618 509782 510854
rect 509866 510618 510102 510854
rect 509546 474938 509782 475174
rect 509866 474938 510102 475174
rect 509546 474618 509782 474854
rect 509866 474618 510102 474854
rect 509546 438938 509782 439174
rect 509866 438938 510102 439174
rect 509546 438618 509782 438854
rect 509866 438618 510102 438854
rect 509546 402938 509782 403174
rect 509866 402938 510102 403174
rect 509546 402618 509782 402854
rect 509866 402618 510102 402854
rect 509546 366938 509782 367174
rect 509866 366938 510102 367174
rect 509546 366618 509782 366854
rect 509866 366618 510102 366854
rect 509546 330938 509782 331174
rect 509866 330938 510102 331174
rect 509546 330618 509782 330854
rect 509866 330618 510102 330854
rect 509546 294938 509782 295174
rect 509866 294938 510102 295174
rect 509546 294618 509782 294854
rect 509866 294618 510102 294854
rect 509546 258938 509782 259174
rect 509866 258938 510102 259174
rect 509546 258618 509782 258854
rect 509866 258618 510102 258854
rect 509546 222938 509782 223174
rect 509866 222938 510102 223174
rect 509546 222618 509782 222854
rect 509866 222618 510102 222854
rect 509546 186938 509782 187174
rect 509866 186938 510102 187174
rect 509546 186618 509782 186854
rect 509866 186618 510102 186854
rect 509546 150938 509782 151174
rect 509866 150938 510102 151174
rect 509546 150618 509782 150854
rect 509866 150618 510102 150854
rect 509546 114938 509782 115174
rect 509866 114938 510102 115174
rect 509546 114618 509782 114854
rect 509866 114618 510102 114854
rect 509546 78938 509782 79174
rect 509866 78938 510102 79174
rect 509546 78618 509782 78854
rect 509866 78618 510102 78854
rect 509546 42938 509782 43174
rect 509866 42938 510102 43174
rect 509546 42618 509782 42854
rect 509866 42618 510102 42854
rect 509546 6938 509782 7174
rect 509866 6938 510102 7174
rect 509546 6618 509782 6854
rect 509866 6618 510102 6854
rect 509546 -2502 509782 -2266
rect 509866 -2502 510102 -2266
rect 509546 -2822 509782 -2586
rect 509866 -2822 510102 -2586
rect 513266 694658 513502 694894
rect 513586 694658 513822 694894
rect 513266 694338 513502 694574
rect 513586 694338 513822 694574
rect 513266 658658 513502 658894
rect 513586 658658 513822 658894
rect 513266 658338 513502 658574
rect 513586 658338 513822 658574
rect 513266 622658 513502 622894
rect 513586 622658 513822 622894
rect 513266 622338 513502 622574
rect 513586 622338 513822 622574
rect 513266 586658 513502 586894
rect 513586 586658 513822 586894
rect 513266 586338 513502 586574
rect 513586 586338 513822 586574
rect 513266 550658 513502 550894
rect 513586 550658 513822 550894
rect 513266 550338 513502 550574
rect 513586 550338 513822 550574
rect 513266 514658 513502 514894
rect 513586 514658 513822 514894
rect 513266 514338 513502 514574
rect 513586 514338 513822 514574
rect 513266 478658 513502 478894
rect 513586 478658 513822 478894
rect 513266 478338 513502 478574
rect 513586 478338 513822 478574
rect 513266 442658 513502 442894
rect 513586 442658 513822 442894
rect 513266 442338 513502 442574
rect 513586 442338 513822 442574
rect 513266 406658 513502 406894
rect 513586 406658 513822 406894
rect 513266 406338 513502 406574
rect 513586 406338 513822 406574
rect 513266 370658 513502 370894
rect 513586 370658 513822 370894
rect 513266 370338 513502 370574
rect 513586 370338 513822 370574
rect 513266 334658 513502 334894
rect 513586 334658 513822 334894
rect 513266 334338 513502 334574
rect 513586 334338 513822 334574
rect 513266 298658 513502 298894
rect 513586 298658 513822 298894
rect 513266 298338 513502 298574
rect 513586 298338 513822 298574
rect 513266 262658 513502 262894
rect 513586 262658 513822 262894
rect 513266 262338 513502 262574
rect 513586 262338 513822 262574
rect 513266 226658 513502 226894
rect 513586 226658 513822 226894
rect 513266 226338 513502 226574
rect 513586 226338 513822 226574
rect 513266 190658 513502 190894
rect 513586 190658 513822 190894
rect 513266 190338 513502 190574
rect 513586 190338 513822 190574
rect 513266 154658 513502 154894
rect 513586 154658 513822 154894
rect 513266 154338 513502 154574
rect 513586 154338 513822 154574
rect 513266 118658 513502 118894
rect 513586 118658 513822 118894
rect 513266 118338 513502 118574
rect 513586 118338 513822 118574
rect 513266 82658 513502 82894
rect 513586 82658 513822 82894
rect 513266 82338 513502 82574
rect 513586 82338 513822 82574
rect 513266 46658 513502 46894
rect 513586 46658 513822 46894
rect 513266 46338 513502 46574
rect 513586 46338 513822 46574
rect 513266 10658 513502 10894
rect 513586 10658 513822 10894
rect 513266 10338 513502 10574
rect 513586 10338 513822 10574
rect 513266 -4422 513502 -4186
rect 513586 -4422 513822 -4186
rect 513266 -4742 513502 -4506
rect 513586 -4742 513822 -4506
rect 534986 711322 535222 711558
rect 535306 711322 535542 711558
rect 534986 711002 535222 711238
rect 535306 711002 535542 711238
rect 531266 709402 531502 709638
rect 531586 709402 531822 709638
rect 531266 709082 531502 709318
rect 531586 709082 531822 709318
rect 527546 707482 527782 707718
rect 527866 707482 528102 707718
rect 527546 707162 527782 707398
rect 527866 707162 528102 707398
rect 516986 698378 517222 698614
rect 517306 698378 517542 698614
rect 516986 698058 517222 698294
rect 517306 698058 517542 698294
rect 516986 662378 517222 662614
rect 517306 662378 517542 662614
rect 516986 662058 517222 662294
rect 517306 662058 517542 662294
rect 516986 626378 517222 626614
rect 517306 626378 517542 626614
rect 516986 626058 517222 626294
rect 517306 626058 517542 626294
rect 516986 590378 517222 590614
rect 517306 590378 517542 590614
rect 516986 590058 517222 590294
rect 517306 590058 517542 590294
rect 516986 554378 517222 554614
rect 517306 554378 517542 554614
rect 516986 554058 517222 554294
rect 517306 554058 517542 554294
rect 516986 518378 517222 518614
rect 517306 518378 517542 518614
rect 516986 518058 517222 518294
rect 517306 518058 517542 518294
rect 516986 482378 517222 482614
rect 517306 482378 517542 482614
rect 516986 482058 517222 482294
rect 517306 482058 517542 482294
rect 516986 446378 517222 446614
rect 517306 446378 517542 446614
rect 516986 446058 517222 446294
rect 517306 446058 517542 446294
rect 516986 410378 517222 410614
rect 517306 410378 517542 410614
rect 516986 410058 517222 410294
rect 517306 410058 517542 410294
rect 516986 374378 517222 374614
rect 517306 374378 517542 374614
rect 516986 374058 517222 374294
rect 517306 374058 517542 374294
rect 516986 338378 517222 338614
rect 517306 338378 517542 338614
rect 516986 338058 517222 338294
rect 517306 338058 517542 338294
rect 516986 302378 517222 302614
rect 517306 302378 517542 302614
rect 516986 302058 517222 302294
rect 517306 302058 517542 302294
rect 516986 266378 517222 266614
rect 517306 266378 517542 266614
rect 516986 266058 517222 266294
rect 517306 266058 517542 266294
rect 516986 230378 517222 230614
rect 517306 230378 517542 230614
rect 516986 230058 517222 230294
rect 517306 230058 517542 230294
rect 516986 194378 517222 194614
rect 517306 194378 517542 194614
rect 516986 194058 517222 194294
rect 517306 194058 517542 194294
rect 516986 158378 517222 158614
rect 517306 158378 517542 158614
rect 516986 158058 517222 158294
rect 517306 158058 517542 158294
rect 516986 122378 517222 122614
rect 517306 122378 517542 122614
rect 516986 122058 517222 122294
rect 517306 122058 517542 122294
rect 516986 86378 517222 86614
rect 517306 86378 517542 86614
rect 516986 86058 517222 86294
rect 517306 86058 517542 86294
rect 516986 50378 517222 50614
rect 517306 50378 517542 50614
rect 516986 50058 517222 50294
rect 517306 50058 517542 50294
rect 516986 14378 517222 14614
rect 517306 14378 517542 14614
rect 516986 14058 517222 14294
rect 517306 14058 517542 14294
rect 498986 -7302 499222 -7066
rect 499306 -7302 499542 -7066
rect 498986 -7622 499222 -7386
rect 499306 -7622 499542 -7386
rect 523826 705562 524062 705798
rect 524146 705562 524382 705798
rect 523826 705242 524062 705478
rect 524146 705242 524382 705478
rect 523826 669218 524062 669454
rect 524146 669218 524382 669454
rect 523826 668898 524062 669134
rect 524146 668898 524382 669134
rect 523826 633218 524062 633454
rect 524146 633218 524382 633454
rect 523826 632898 524062 633134
rect 524146 632898 524382 633134
rect 523826 597218 524062 597454
rect 524146 597218 524382 597454
rect 523826 596898 524062 597134
rect 524146 596898 524382 597134
rect 523826 561218 524062 561454
rect 524146 561218 524382 561454
rect 523826 560898 524062 561134
rect 524146 560898 524382 561134
rect 523826 525218 524062 525454
rect 524146 525218 524382 525454
rect 523826 524898 524062 525134
rect 524146 524898 524382 525134
rect 523826 489218 524062 489454
rect 524146 489218 524382 489454
rect 523826 488898 524062 489134
rect 524146 488898 524382 489134
rect 523826 453218 524062 453454
rect 524146 453218 524382 453454
rect 523826 452898 524062 453134
rect 524146 452898 524382 453134
rect 523826 417218 524062 417454
rect 524146 417218 524382 417454
rect 523826 416898 524062 417134
rect 524146 416898 524382 417134
rect 523826 381218 524062 381454
rect 524146 381218 524382 381454
rect 523826 380898 524062 381134
rect 524146 380898 524382 381134
rect 523826 345218 524062 345454
rect 524146 345218 524382 345454
rect 523826 344898 524062 345134
rect 524146 344898 524382 345134
rect 523826 309218 524062 309454
rect 524146 309218 524382 309454
rect 523826 308898 524062 309134
rect 524146 308898 524382 309134
rect 523826 273218 524062 273454
rect 524146 273218 524382 273454
rect 523826 272898 524062 273134
rect 524146 272898 524382 273134
rect 523826 237218 524062 237454
rect 524146 237218 524382 237454
rect 523826 236898 524062 237134
rect 524146 236898 524382 237134
rect 523826 201218 524062 201454
rect 524146 201218 524382 201454
rect 523826 200898 524062 201134
rect 524146 200898 524382 201134
rect 523826 165218 524062 165454
rect 524146 165218 524382 165454
rect 523826 164898 524062 165134
rect 524146 164898 524382 165134
rect 523826 129218 524062 129454
rect 524146 129218 524382 129454
rect 523826 128898 524062 129134
rect 524146 128898 524382 129134
rect 523826 93218 524062 93454
rect 524146 93218 524382 93454
rect 523826 92898 524062 93134
rect 524146 92898 524382 93134
rect 523826 57218 524062 57454
rect 524146 57218 524382 57454
rect 523826 56898 524062 57134
rect 524146 56898 524382 57134
rect 523826 21218 524062 21454
rect 524146 21218 524382 21454
rect 523826 20898 524062 21134
rect 524146 20898 524382 21134
rect 523826 -1542 524062 -1306
rect 524146 -1542 524382 -1306
rect 523826 -1862 524062 -1626
rect 524146 -1862 524382 -1626
rect 527546 672938 527782 673174
rect 527866 672938 528102 673174
rect 527546 672618 527782 672854
rect 527866 672618 528102 672854
rect 527546 636938 527782 637174
rect 527866 636938 528102 637174
rect 527546 636618 527782 636854
rect 527866 636618 528102 636854
rect 527546 600938 527782 601174
rect 527866 600938 528102 601174
rect 527546 600618 527782 600854
rect 527866 600618 528102 600854
rect 527546 564938 527782 565174
rect 527866 564938 528102 565174
rect 527546 564618 527782 564854
rect 527866 564618 528102 564854
rect 527546 528938 527782 529174
rect 527866 528938 528102 529174
rect 527546 528618 527782 528854
rect 527866 528618 528102 528854
rect 527546 492938 527782 493174
rect 527866 492938 528102 493174
rect 527546 492618 527782 492854
rect 527866 492618 528102 492854
rect 527546 456938 527782 457174
rect 527866 456938 528102 457174
rect 527546 456618 527782 456854
rect 527866 456618 528102 456854
rect 527546 420938 527782 421174
rect 527866 420938 528102 421174
rect 527546 420618 527782 420854
rect 527866 420618 528102 420854
rect 527546 384938 527782 385174
rect 527866 384938 528102 385174
rect 527546 384618 527782 384854
rect 527866 384618 528102 384854
rect 527546 348938 527782 349174
rect 527866 348938 528102 349174
rect 527546 348618 527782 348854
rect 527866 348618 528102 348854
rect 527546 312938 527782 313174
rect 527866 312938 528102 313174
rect 527546 312618 527782 312854
rect 527866 312618 528102 312854
rect 527546 276938 527782 277174
rect 527866 276938 528102 277174
rect 527546 276618 527782 276854
rect 527866 276618 528102 276854
rect 527546 240938 527782 241174
rect 527866 240938 528102 241174
rect 527546 240618 527782 240854
rect 527866 240618 528102 240854
rect 527546 204938 527782 205174
rect 527866 204938 528102 205174
rect 527546 204618 527782 204854
rect 527866 204618 528102 204854
rect 527546 168938 527782 169174
rect 527866 168938 528102 169174
rect 527546 168618 527782 168854
rect 527866 168618 528102 168854
rect 527546 132938 527782 133174
rect 527866 132938 528102 133174
rect 527546 132618 527782 132854
rect 527866 132618 528102 132854
rect 527546 96938 527782 97174
rect 527866 96938 528102 97174
rect 527546 96618 527782 96854
rect 527866 96618 528102 96854
rect 527546 60938 527782 61174
rect 527866 60938 528102 61174
rect 527546 60618 527782 60854
rect 527866 60618 528102 60854
rect 527546 24938 527782 25174
rect 527866 24938 528102 25174
rect 527546 24618 527782 24854
rect 527866 24618 528102 24854
rect 527546 -3462 527782 -3226
rect 527866 -3462 528102 -3226
rect 527546 -3782 527782 -3546
rect 527866 -3782 528102 -3546
rect 531266 676658 531502 676894
rect 531586 676658 531822 676894
rect 531266 676338 531502 676574
rect 531586 676338 531822 676574
rect 531266 640658 531502 640894
rect 531586 640658 531822 640894
rect 531266 640338 531502 640574
rect 531586 640338 531822 640574
rect 531266 604658 531502 604894
rect 531586 604658 531822 604894
rect 531266 604338 531502 604574
rect 531586 604338 531822 604574
rect 531266 568658 531502 568894
rect 531586 568658 531822 568894
rect 531266 568338 531502 568574
rect 531586 568338 531822 568574
rect 531266 532658 531502 532894
rect 531586 532658 531822 532894
rect 531266 532338 531502 532574
rect 531586 532338 531822 532574
rect 531266 496658 531502 496894
rect 531586 496658 531822 496894
rect 531266 496338 531502 496574
rect 531586 496338 531822 496574
rect 531266 460658 531502 460894
rect 531586 460658 531822 460894
rect 531266 460338 531502 460574
rect 531586 460338 531822 460574
rect 531266 424658 531502 424894
rect 531586 424658 531822 424894
rect 531266 424338 531502 424574
rect 531586 424338 531822 424574
rect 531266 388658 531502 388894
rect 531586 388658 531822 388894
rect 531266 388338 531502 388574
rect 531586 388338 531822 388574
rect 531266 352658 531502 352894
rect 531586 352658 531822 352894
rect 531266 352338 531502 352574
rect 531586 352338 531822 352574
rect 531266 316658 531502 316894
rect 531586 316658 531822 316894
rect 531266 316338 531502 316574
rect 531586 316338 531822 316574
rect 531266 280658 531502 280894
rect 531586 280658 531822 280894
rect 531266 280338 531502 280574
rect 531586 280338 531822 280574
rect 531266 244658 531502 244894
rect 531586 244658 531822 244894
rect 531266 244338 531502 244574
rect 531586 244338 531822 244574
rect 531266 208658 531502 208894
rect 531586 208658 531822 208894
rect 531266 208338 531502 208574
rect 531586 208338 531822 208574
rect 531266 172658 531502 172894
rect 531586 172658 531822 172894
rect 531266 172338 531502 172574
rect 531586 172338 531822 172574
rect 531266 136658 531502 136894
rect 531586 136658 531822 136894
rect 531266 136338 531502 136574
rect 531586 136338 531822 136574
rect 531266 100658 531502 100894
rect 531586 100658 531822 100894
rect 531266 100338 531502 100574
rect 531586 100338 531822 100574
rect 531266 64658 531502 64894
rect 531586 64658 531822 64894
rect 531266 64338 531502 64574
rect 531586 64338 531822 64574
rect 531266 28658 531502 28894
rect 531586 28658 531822 28894
rect 531266 28338 531502 28574
rect 531586 28338 531822 28574
rect 531266 -5382 531502 -5146
rect 531586 -5382 531822 -5146
rect 531266 -5702 531502 -5466
rect 531586 -5702 531822 -5466
rect 552986 710362 553222 710598
rect 553306 710362 553542 710598
rect 552986 710042 553222 710278
rect 553306 710042 553542 710278
rect 549266 708442 549502 708678
rect 549586 708442 549822 708678
rect 549266 708122 549502 708358
rect 549586 708122 549822 708358
rect 545546 706522 545782 706758
rect 545866 706522 546102 706758
rect 545546 706202 545782 706438
rect 545866 706202 546102 706438
rect 534986 680378 535222 680614
rect 535306 680378 535542 680614
rect 534986 680058 535222 680294
rect 535306 680058 535542 680294
rect 534986 644378 535222 644614
rect 535306 644378 535542 644614
rect 534986 644058 535222 644294
rect 535306 644058 535542 644294
rect 534986 608378 535222 608614
rect 535306 608378 535542 608614
rect 534986 608058 535222 608294
rect 535306 608058 535542 608294
rect 534986 572378 535222 572614
rect 535306 572378 535542 572614
rect 534986 572058 535222 572294
rect 535306 572058 535542 572294
rect 534986 536378 535222 536614
rect 535306 536378 535542 536614
rect 534986 536058 535222 536294
rect 535306 536058 535542 536294
rect 534986 500378 535222 500614
rect 535306 500378 535542 500614
rect 534986 500058 535222 500294
rect 535306 500058 535542 500294
rect 534986 464378 535222 464614
rect 535306 464378 535542 464614
rect 534986 464058 535222 464294
rect 535306 464058 535542 464294
rect 534986 428378 535222 428614
rect 535306 428378 535542 428614
rect 534986 428058 535222 428294
rect 535306 428058 535542 428294
rect 534986 392378 535222 392614
rect 535306 392378 535542 392614
rect 534986 392058 535222 392294
rect 535306 392058 535542 392294
rect 534986 356378 535222 356614
rect 535306 356378 535542 356614
rect 534986 356058 535222 356294
rect 535306 356058 535542 356294
rect 534986 320378 535222 320614
rect 535306 320378 535542 320614
rect 534986 320058 535222 320294
rect 535306 320058 535542 320294
rect 534986 284378 535222 284614
rect 535306 284378 535542 284614
rect 534986 284058 535222 284294
rect 535306 284058 535542 284294
rect 534986 248378 535222 248614
rect 535306 248378 535542 248614
rect 534986 248058 535222 248294
rect 535306 248058 535542 248294
rect 534986 212378 535222 212614
rect 535306 212378 535542 212614
rect 534986 212058 535222 212294
rect 535306 212058 535542 212294
rect 534986 176378 535222 176614
rect 535306 176378 535542 176614
rect 534986 176058 535222 176294
rect 535306 176058 535542 176294
rect 534986 140378 535222 140614
rect 535306 140378 535542 140614
rect 534986 140058 535222 140294
rect 535306 140058 535542 140294
rect 534986 104378 535222 104614
rect 535306 104378 535542 104614
rect 534986 104058 535222 104294
rect 535306 104058 535542 104294
rect 534986 68378 535222 68614
rect 535306 68378 535542 68614
rect 534986 68058 535222 68294
rect 535306 68058 535542 68294
rect 534986 32378 535222 32614
rect 535306 32378 535542 32614
rect 534986 32058 535222 32294
rect 535306 32058 535542 32294
rect 516986 -6342 517222 -6106
rect 517306 -6342 517542 -6106
rect 516986 -6662 517222 -6426
rect 517306 -6662 517542 -6426
rect 541826 704602 542062 704838
rect 542146 704602 542382 704838
rect 541826 704282 542062 704518
rect 542146 704282 542382 704518
rect 541826 687218 542062 687454
rect 542146 687218 542382 687454
rect 541826 686898 542062 687134
rect 542146 686898 542382 687134
rect 541826 651218 542062 651454
rect 542146 651218 542382 651454
rect 541826 650898 542062 651134
rect 542146 650898 542382 651134
rect 541826 615218 542062 615454
rect 542146 615218 542382 615454
rect 541826 614898 542062 615134
rect 542146 614898 542382 615134
rect 541826 579218 542062 579454
rect 542146 579218 542382 579454
rect 541826 578898 542062 579134
rect 542146 578898 542382 579134
rect 541826 543218 542062 543454
rect 542146 543218 542382 543454
rect 541826 542898 542062 543134
rect 542146 542898 542382 543134
rect 541826 507218 542062 507454
rect 542146 507218 542382 507454
rect 541826 506898 542062 507134
rect 542146 506898 542382 507134
rect 541826 471218 542062 471454
rect 542146 471218 542382 471454
rect 541826 470898 542062 471134
rect 542146 470898 542382 471134
rect 541826 435218 542062 435454
rect 542146 435218 542382 435454
rect 541826 434898 542062 435134
rect 542146 434898 542382 435134
rect 541826 399218 542062 399454
rect 542146 399218 542382 399454
rect 541826 398898 542062 399134
rect 542146 398898 542382 399134
rect 541826 363218 542062 363454
rect 542146 363218 542382 363454
rect 541826 362898 542062 363134
rect 542146 362898 542382 363134
rect 541826 327218 542062 327454
rect 542146 327218 542382 327454
rect 541826 326898 542062 327134
rect 542146 326898 542382 327134
rect 541826 291218 542062 291454
rect 542146 291218 542382 291454
rect 541826 290898 542062 291134
rect 542146 290898 542382 291134
rect 541826 255218 542062 255454
rect 542146 255218 542382 255454
rect 541826 254898 542062 255134
rect 542146 254898 542382 255134
rect 541826 219218 542062 219454
rect 542146 219218 542382 219454
rect 541826 218898 542062 219134
rect 542146 218898 542382 219134
rect 541826 183218 542062 183454
rect 542146 183218 542382 183454
rect 541826 182898 542062 183134
rect 542146 182898 542382 183134
rect 541826 147218 542062 147454
rect 542146 147218 542382 147454
rect 541826 146898 542062 147134
rect 542146 146898 542382 147134
rect 541826 111218 542062 111454
rect 542146 111218 542382 111454
rect 541826 110898 542062 111134
rect 542146 110898 542382 111134
rect 541826 75218 542062 75454
rect 542146 75218 542382 75454
rect 541826 74898 542062 75134
rect 542146 74898 542382 75134
rect 541826 39218 542062 39454
rect 542146 39218 542382 39454
rect 541826 38898 542062 39134
rect 542146 38898 542382 39134
rect 541826 3218 542062 3454
rect 542146 3218 542382 3454
rect 541826 2898 542062 3134
rect 542146 2898 542382 3134
rect 541826 -582 542062 -346
rect 542146 -582 542382 -346
rect 541826 -902 542062 -666
rect 542146 -902 542382 -666
rect 545546 690938 545782 691174
rect 545866 690938 546102 691174
rect 545546 690618 545782 690854
rect 545866 690618 546102 690854
rect 545546 654938 545782 655174
rect 545866 654938 546102 655174
rect 545546 654618 545782 654854
rect 545866 654618 546102 654854
rect 545546 618938 545782 619174
rect 545866 618938 546102 619174
rect 545546 618618 545782 618854
rect 545866 618618 546102 618854
rect 545546 582938 545782 583174
rect 545866 582938 546102 583174
rect 545546 582618 545782 582854
rect 545866 582618 546102 582854
rect 545546 546938 545782 547174
rect 545866 546938 546102 547174
rect 545546 546618 545782 546854
rect 545866 546618 546102 546854
rect 545546 510938 545782 511174
rect 545866 510938 546102 511174
rect 545546 510618 545782 510854
rect 545866 510618 546102 510854
rect 545546 474938 545782 475174
rect 545866 474938 546102 475174
rect 545546 474618 545782 474854
rect 545866 474618 546102 474854
rect 545546 438938 545782 439174
rect 545866 438938 546102 439174
rect 545546 438618 545782 438854
rect 545866 438618 546102 438854
rect 545546 402938 545782 403174
rect 545866 402938 546102 403174
rect 545546 402618 545782 402854
rect 545866 402618 546102 402854
rect 545546 366938 545782 367174
rect 545866 366938 546102 367174
rect 545546 366618 545782 366854
rect 545866 366618 546102 366854
rect 545546 330938 545782 331174
rect 545866 330938 546102 331174
rect 545546 330618 545782 330854
rect 545866 330618 546102 330854
rect 545546 294938 545782 295174
rect 545866 294938 546102 295174
rect 545546 294618 545782 294854
rect 545866 294618 546102 294854
rect 545546 258938 545782 259174
rect 545866 258938 546102 259174
rect 545546 258618 545782 258854
rect 545866 258618 546102 258854
rect 545546 222938 545782 223174
rect 545866 222938 546102 223174
rect 545546 222618 545782 222854
rect 545866 222618 546102 222854
rect 545546 186938 545782 187174
rect 545866 186938 546102 187174
rect 545546 186618 545782 186854
rect 545866 186618 546102 186854
rect 545546 150938 545782 151174
rect 545866 150938 546102 151174
rect 545546 150618 545782 150854
rect 545866 150618 546102 150854
rect 545546 114938 545782 115174
rect 545866 114938 546102 115174
rect 545546 114618 545782 114854
rect 545866 114618 546102 114854
rect 545546 78938 545782 79174
rect 545866 78938 546102 79174
rect 545546 78618 545782 78854
rect 545866 78618 546102 78854
rect 545546 42938 545782 43174
rect 545866 42938 546102 43174
rect 545546 42618 545782 42854
rect 545866 42618 546102 42854
rect 545546 6938 545782 7174
rect 545866 6938 546102 7174
rect 545546 6618 545782 6854
rect 545866 6618 546102 6854
rect 545546 -2502 545782 -2266
rect 545866 -2502 546102 -2266
rect 545546 -2822 545782 -2586
rect 545866 -2822 546102 -2586
rect 549266 694658 549502 694894
rect 549586 694658 549822 694894
rect 549266 694338 549502 694574
rect 549586 694338 549822 694574
rect 549266 658658 549502 658894
rect 549586 658658 549822 658894
rect 549266 658338 549502 658574
rect 549586 658338 549822 658574
rect 549266 622658 549502 622894
rect 549586 622658 549822 622894
rect 549266 622338 549502 622574
rect 549586 622338 549822 622574
rect 549266 586658 549502 586894
rect 549586 586658 549822 586894
rect 549266 586338 549502 586574
rect 549586 586338 549822 586574
rect 549266 550658 549502 550894
rect 549586 550658 549822 550894
rect 549266 550338 549502 550574
rect 549586 550338 549822 550574
rect 549266 514658 549502 514894
rect 549586 514658 549822 514894
rect 549266 514338 549502 514574
rect 549586 514338 549822 514574
rect 549266 478658 549502 478894
rect 549586 478658 549822 478894
rect 549266 478338 549502 478574
rect 549586 478338 549822 478574
rect 549266 442658 549502 442894
rect 549586 442658 549822 442894
rect 549266 442338 549502 442574
rect 549586 442338 549822 442574
rect 549266 406658 549502 406894
rect 549586 406658 549822 406894
rect 549266 406338 549502 406574
rect 549586 406338 549822 406574
rect 549266 370658 549502 370894
rect 549586 370658 549822 370894
rect 549266 370338 549502 370574
rect 549586 370338 549822 370574
rect 549266 334658 549502 334894
rect 549586 334658 549822 334894
rect 549266 334338 549502 334574
rect 549586 334338 549822 334574
rect 549266 298658 549502 298894
rect 549586 298658 549822 298894
rect 549266 298338 549502 298574
rect 549586 298338 549822 298574
rect 549266 262658 549502 262894
rect 549586 262658 549822 262894
rect 549266 262338 549502 262574
rect 549586 262338 549822 262574
rect 549266 226658 549502 226894
rect 549586 226658 549822 226894
rect 549266 226338 549502 226574
rect 549586 226338 549822 226574
rect 549266 190658 549502 190894
rect 549586 190658 549822 190894
rect 549266 190338 549502 190574
rect 549586 190338 549822 190574
rect 549266 154658 549502 154894
rect 549586 154658 549822 154894
rect 549266 154338 549502 154574
rect 549586 154338 549822 154574
rect 549266 118658 549502 118894
rect 549586 118658 549822 118894
rect 549266 118338 549502 118574
rect 549586 118338 549822 118574
rect 549266 82658 549502 82894
rect 549586 82658 549822 82894
rect 549266 82338 549502 82574
rect 549586 82338 549822 82574
rect 549266 46658 549502 46894
rect 549586 46658 549822 46894
rect 549266 46338 549502 46574
rect 549586 46338 549822 46574
rect 549266 10658 549502 10894
rect 549586 10658 549822 10894
rect 549266 10338 549502 10574
rect 549586 10338 549822 10574
rect 549266 -4422 549502 -4186
rect 549586 -4422 549822 -4186
rect 549266 -4742 549502 -4506
rect 549586 -4742 549822 -4506
rect 570986 711322 571222 711558
rect 571306 711322 571542 711558
rect 570986 711002 571222 711238
rect 571306 711002 571542 711238
rect 567266 709402 567502 709638
rect 567586 709402 567822 709638
rect 567266 709082 567502 709318
rect 567586 709082 567822 709318
rect 563546 707482 563782 707718
rect 563866 707482 564102 707718
rect 563546 707162 563782 707398
rect 563866 707162 564102 707398
rect 552986 698378 553222 698614
rect 553306 698378 553542 698614
rect 552986 698058 553222 698294
rect 553306 698058 553542 698294
rect 552986 662378 553222 662614
rect 553306 662378 553542 662614
rect 552986 662058 553222 662294
rect 553306 662058 553542 662294
rect 552986 626378 553222 626614
rect 553306 626378 553542 626614
rect 552986 626058 553222 626294
rect 553306 626058 553542 626294
rect 552986 590378 553222 590614
rect 553306 590378 553542 590614
rect 552986 590058 553222 590294
rect 553306 590058 553542 590294
rect 552986 554378 553222 554614
rect 553306 554378 553542 554614
rect 552986 554058 553222 554294
rect 553306 554058 553542 554294
rect 552986 518378 553222 518614
rect 553306 518378 553542 518614
rect 552986 518058 553222 518294
rect 553306 518058 553542 518294
rect 552986 482378 553222 482614
rect 553306 482378 553542 482614
rect 552986 482058 553222 482294
rect 553306 482058 553542 482294
rect 552986 446378 553222 446614
rect 553306 446378 553542 446614
rect 552986 446058 553222 446294
rect 553306 446058 553542 446294
rect 552986 410378 553222 410614
rect 553306 410378 553542 410614
rect 552986 410058 553222 410294
rect 553306 410058 553542 410294
rect 552986 374378 553222 374614
rect 553306 374378 553542 374614
rect 552986 374058 553222 374294
rect 553306 374058 553542 374294
rect 552986 338378 553222 338614
rect 553306 338378 553542 338614
rect 552986 338058 553222 338294
rect 553306 338058 553542 338294
rect 552986 302378 553222 302614
rect 553306 302378 553542 302614
rect 552986 302058 553222 302294
rect 553306 302058 553542 302294
rect 552986 266378 553222 266614
rect 553306 266378 553542 266614
rect 552986 266058 553222 266294
rect 553306 266058 553542 266294
rect 552986 230378 553222 230614
rect 553306 230378 553542 230614
rect 552986 230058 553222 230294
rect 553306 230058 553542 230294
rect 552986 194378 553222 194614
rect 553306 194378 553542 194614
rect 552986 194058 553222 194294
rect 553306 194058 553542 194294
rect 552986 158378 553222 158614
rect 553306 158378 553542 158614
rect 552986 158058 553222 158294
rect 553306 158058 553542 158294
rect 552986 122378 553222 122614
rect 553306 122378 553542 122614
rect 552986 122058 553222 122294
rect 553306 122058 553542 122294
rect 552986 86378 553222 86614
rect 553306 86378 553542 86614
rect 552986 86058 553222 86294
rect 553306 86058 553542 86294
rect 552986 50378 553222 50614
rect 553306 50378 553542 50614
rect 552986 50058 553222 50294
rect 553306 50058 553542 50294
rect 552986 14378 553222 14614
rect 553306 14378 553542 14614
rect 552986 14058 553222 14294
rect 553306 14058 553542 14294
rect 534986 -7302 535222 -7066
rect 535306 -7302 535542 -7066
rect 534986 -7622 535222 -7386
rect 535306 -7622 535542 -7386
rect 559826 705562 560062 705798
rect 560146 705562 560382 705798
rect 559826 705242 560062 705478
rect 560146 705242 560382 705478
rect 559826 669218 560062 669454
rect 560146 669218 560382 669454
rect 559826 668898 560062 669134
rect 560146 668898 560382 669134
rect 559826 633218 560062 633454
rect 560146 633218 560382 633454
rect 559826 632898 560062 633134
rect 560146 632898 560382 633134
rect 559826 597218 560062 597454
rect 560146 597218 560382 597454
rect 559826 596898 560062 597134
rect 560146 596898 560382 597134
rect 559826 561218 560062 561454
rect 560146 561218 560382 561454
rect 559826 560898 560062 561134
rect 560146 560898 560382 561134
rect 559826 525218 560062 525454
rect 560146 525218 560382 525454
rect 559826 524898 560062 525134
rect 560146 524898 560382 525134
rect 559826 489218 560062 489454
rect 560146 489218 560382 489454
rect 559826 488898 560062 489134
rect 560146 488898 560382 489134
rect 559826 453218 560062 453454
rect 560146 453218 560382 453454
rect 559826 452898 560062 453134
rect 560146 452898 560382 453134
rect 559826 417218 560062 417454
rect 560146 417218 560382 417454
rect 559826 416898 560062 417134
rect 560146 416898 560382 417134
rect 559826 381218 560062 381454
rect 560146 381218 560382 381454
rect 559826 380898 560062 381134
rect 560146 380898 560382 381134
rect 559826 345218 560062 345454
rect 560146 345218 560382 345454
rect 559826 344898 560062 345134
rect 560146 344898 560382 345134
rect 559826 309218 560062 309454
rect 560146 309218 560382 309454
rect 559826 308898 560062 309134
rect 560146 308898 560382 309134
rect 559826 273218 560062 273454
rect 560146 273218 560382 273454
rect 559826 272898 560062 273134
rect 560146 272898 560382 273134
rect 559826 237218 560062 237454
rect 560146 237218 560382 237454
rect 559826 236898 560062 237134
rect 560146 236898 560382 237134
rect 559826 201218 560062 201454
rect 560146 201218 560382 201454
rect 559826 200898 560062 201134
rect 560146 200898 560382 201134
rect 559826 165218 560062 165454
rect 560146 165218 560382 165454
rect 559826 164898 560062 165134
rect 560146 164898 560382 165134
rect 559826 129218 560062 129454
rect 560146 129218 560382 129454
rect 559826 128898 560062 129134
rect 560146 128898 560382 129134
rect 559826 93218 560062 93454
rect 560146 93218 560382 93454
rect 559826 92898 560062 93134
rect 560146 92898 560382 93134
rect 559826 57218 560062 57454
rect 560146 57218 560382 57454
rect 559826 56898 560062 57134
rect 560146 56898 560382 57134
rect 559826 21218 560062 21454
rect 560146 21218 560382 21454
rect 559826 20898 560062 21134
rect 560146 20898 560382 21134
rect 559826 -1542 560062 -1306
rect 560146 -1542 560382 -1306
rect 559826 -1862 560062 -1626
rect 560146 -1862 560382 -1626
rect 563546 672938 563782 673174
rect 563866 672938 564102 673174
rect 563546 672618 563782 672854
rect 563866 672618 564102 672854
rect 563546 636938 563782 637174
rect 563866 636938 564102 637174
rect 563546 636618 563782 636854
rect 563866 636618 564102 636854
rect 563546 600938 563782 601174
rect 563866 600938 564102 601174
rect 563546 600618 563782 600854
rect 563866 600618 564102 600854
rect 563546 564938 563782 565174
rect 563866 564938 564102 565174
rect 563546 564618 563782 564854
rect 563866 564618 564102 564854
rect 563546 528938 563782 529174
rect 563866 528938 564102 529174
rect 563546 528618 563782 528854
rect 563866 528618 564102 528854
rect 563546 492938 563782 493174
rect 563866 492938 564102 493174
rect 563546 492618 563782 492854
rect 563866 492618 564102 492854
rect 563546 456938 563782 457174
rect 563866 456938 564102 457174
rect 563546 456618 563782 456854
rect 563866 456618 564102 456854
rect 563546 420938 563782 421174
rect 563866 420938 564102 421174
rect 563546 420618 563782 420854
rect 563866 420618 564102 420854
rect 563546 384938 563782 385174
rect 563866 384938 564102 385174
rect 563546 384618 563782 384854
rect 563866 384618 564102 384854
rect 563546 348938 563782 349174
rect 563866 348938 564102 349174
rect 563546 348618 563782 348854
rect 563866 348618 564102 348854
rect 563546 312938 563782 313174
rect 563866 312938 564102 313174
rect 563546 312618 563782 312854
rect 563866 312618 564102 312854
rect 563546 276938 563782 277174
rect 563866 276938 564102 277174
rect 563546 276618 563782 276854
rect 563866 276618 564102 276854
rect 563546 240938 563782 241174
rect 563866 240938 564102 241174
rect 563546 240618 563782 240854
rect 563866 240618 564102 240854
rect 563546 204938 563782 205174
rect 563866 204938 564102 205174
rect 563546 204618 563782 204854
rect 563866 204618 564102 204854
rect 563546 168938 563782 169174
rect 563866 168938 564102 169174
rect 563546 168618 563782 168854
rect 563866 168618 564102 168854
rect 563546 132938 563782 133174
rect 563866 132938 564102 133174
rect 563546 132618 563782 132854
rect 563866 132618 564102 132854
rect 563546 96938 563782 97174
rect 563866 96938 564102 97174
rect 563546 96618 563782 96854
rect 563866 96618 564102 96854
rect 563546 60938 563782 61174
rect 563866 60938 564102 61174
rect 563546 60618 563782 60854
rect 563866 60618 564102 60854
rect 563546 24938 563782 25174
rect 563866 24938 564102 25174
rect 563546 24618 563782 24854
rect 563866 24618 564102 24854
rect 563546 -3462 563782 -3226
rect 563866 -3462 564102 -3226
rect 563546 -3782 563782 -3546
rect 563866 -3782 564102 -3546
rect 567266 676658 567502 676894
rect 567586 676658 567822 676894
rect 567266 676338 567502 676574
rect 567586 676338 567822 676574
rect 567266 640658 567502 640894
rect 567586 640658 567822 640894
rect 567266 640338 567502 640574
rect 567586 640338 567822 640574
rect 567266 604658 567502 604894
rect 567586 604658 567822 604894
rect 567266 604338 567502 604574
rect 567586 604338 567822 604574
rect 567266 568658 567502 568894
rect 567586 568658 567822 568894
rect 567266 568338 567502 568574
rect 567586 568338 567822 568574
rect 567266 532658 567502 532894
rect 567586 532658 567822 532894
rect 567266 532338 567502 532574
rect 567586 532338 567822 532574
rect 567266 496658 567502 496894
rect 567586 496658 567822 496894
rect 567266 496338 567502 496574
rect 567586 496338 567822 496574
rect 567266 460658 567502 460894
rect 567586 460658 567822 460894
rect 567266 460338 567502 460574
rect 567586 460338 567822 460574
rect 567266 424658 567502 424894
rect 567586 424658 567822 424894
rect 567266 424338 567502 424574
rect 567586 424338 567822 424574
rect 567266 388658 567502 388894
rect 567586 388658 567822 388894
rect 567266 388338 567502 388574
rect 567586 388338 567822 388574
rect 567266 352658 567502 352894
rect 567586 352658 567822 352894
rect 567266 352338 567502 352574
rect 567586 352338 567822 352574
rect 567266 316658 567502 316894
rect 567586 316658 567822 316894
rect 567266 316338 567502 316574
rect 567586 316338 567822 316574
rect 567266 280658 567502 280894
rect 567586 280658 567822 280894
rect 567266 280338 567502 280574
rect 567586 280338 567822 280574
rect 567266 244658 567502 244894
rect 567586 244658 567822 244894
rect 567266 244338 567502 244574
rect 567586 244338 567822 244574
rect 567266 208658 567502 208894
rect 567586 208658 567822 208894
rect 567266 208338 567502 208574
rect 567586 208338 567822 208574
rect 567266 172658 567502 172894
rect 567586 172658 567822 172894
rect 567266 172338 567502 172574
rect 567586 172338 567822 172574
rect 567266 136658 567502 136894
rect 567586 136658 567822 136894
rect 567266 136338 567502 136574
rect 567586 136338 567822 136574
rect 567266 100658 567502 100894
rect 567586 100658 567822 100894
rect 567266 100338 567502 100574
rect 567586 100338 567822 100574
rect 567266 64658 567502 64894
rect 567586 64658 567822 64894
rect 567266 64338 567502 64574
rect 567586 64338 567822 64574
rect 567266 28658 567502 28894
rect 567586 28658 567822 28894
rect 567266 28338 567502 28574
rect 567586 28338 567822 28574
rect 567266 -5382 567502 -5146
rect 567586 -5382 567822 -5146
rect 567266 -5702 567502 -5466
rect 567586 -5702 567822 -5466
rect 592062 711322 592298 711558
rect 592382 711322 592618 711558
rect 592062 711002 592298 711238
rect 592382 711002 592618 711238
rect 591102 710362 591338 710598
rect 591422 710362 591658 710598
rect 591102 710042 591338 710278
rect 591422 710042 591658 710278
rect 590142 709402 590378 709638
rect 590462 709402 590698 709638
rect 590142 709082 590378 709318
rect 590462 709082 590698 709318
rect 589182 708442 589418 708678
rect 589502 708442 589738 708678
rect 589182 708122 589418 708358
rect 589502 708122 589738 708358
rect 588222 707482 588458 707718
rect 588542 707482 588778 707718
rect 588222 707162 588458 707398
rect 588542 707162 588778 707398
rect 581546 706522 581782 706758
rect 581866 706522 582102 706758
rect 581546 706202 581782 706438
rect 581866 706202 582102 706438
rect 570986 680378 571222 680614
rect 571306 680378 571542 680614
rect 570986 680058 571222 680294
rect 571306 680058 571542 680294
rect 570986 644378 571222 644614
rect 571306 644378 571542 644614
rect 570986 644058 571222 644294
rect 571306 644058 571542 644294
rect 570986 608378 571222 608614
rect 571306 608378 571542 608614
rect 570986 608058 571222 608294
rect 571306 608058 571542 608294
rect 570986 572378 571222 572614
rect 571306 572378 571542 572614
rect 570986 572058 571222 572294
rect 571306 572058 571542 572294
rect 570986 536378 571222 536614
rect 571306 536378 571542 536614
rect 570986 536058 571222 536294
rect 571306 536058 571542 536294
rect 570986 500378 571222 500614
rect 571306 500378 571542 500614
rect 570986 500058 571222 500294
rect 571306 500058 571542 500294
rect 570986 464378 571222 464614
rect 571306 464378 571542 464614
rect 570986 464058 571222 464294
rect 571306 464058 571542 464294
rect 570986 428378 571222 428614
rect 571306 428378 571542 428614
rect 570986 428058 571222 428294
rect 571306 428058 571542 428294
rect 570986 392378 571222 392614
rect 571306 392378 571542 392614
rect 570986 392058 571222 392294
rect 571306 392058 571542 392294
rect 570986 356378 571222 356614
rect 571306 356378 571542 356614
rect 570986 356058 571222 356294
rect 571306 356058 571542 356294
rect 570986 320378 571222 320614
rect 571306 320378 571542 320614
rect 570986 320058 571222 320294
rect 571306 320058 571542 320294
rect 570986 284378 571222 284614
rect 571306 284378 571542 284614
rect 570986 284058 571222 284294
rect 571306 284058 571542 284294
rect 570986 248378 571222 248614
rect 571306 248378 571542 248614
rect 570986 248058 571222 248294
rect 571306 248058 571542 248294
rect 570986 212378 571222 212614
rect 571306 212378 571542 212614
rect 570986 212058 571222 212294
rect 571306 212058 571542 212294
rect 570986 176378 571222 176614
rect 571306 176378 571542 176614
rect 570986 176058 571222 176294
rect 571306 176058 571542 176294
rect 570986 140378 571222 140614
rect 571306 140378 571542 140614
rect 570986 140058 571222 140294
rect 571306 140058 571542 140294
rect 570986 104378 571222 104614
rect 571306 104378 571542 104614
rect 570986 104058 571222 104294
rect 571306 104058 571542 104294
rect 570986 68378 571222 68614
rect 571306 68378 571542 68614
rect 570986 68058 571222 68294
rect 571306 68058 571542 68294
rect 570986 32378 571222 32614
rect 571306 32378 571542 32614
rect 570986 32058 571222 32294
rect 571306 32058 571542 32294
rect 552986 -6342 553222 -6106
rect 553306 -6342 553542 -6106
rect 552986 -6662 553222 -6426
rect 553306 -6662 553542 -6426
rect 577826 704602 578062 704838
rect 578146 704602 578382 704838
rect 577826 704282 578062 704518
rect 578146 704282 578382 704518
rect 577826 687218 578062 687454
rect 578146 687218 578382 687454
rect 577826 686898 578062 687134
rect 578146 686898 578382 687134
rect 577826 651218 578062 651454
rect 578146 651218 578382 651454
rect 577826 650898 578062 651134
rect 578146 650898 578382 651134
rect 577826 615218 578062 615454
rect 578146 615218 578382 615454
rect 577826 614898 578062 615134
rect 578146 614898 578382 615134
rect 577826 579218 578062 579454
rect 578146 579218 578382 579454
rect 577826 578898 578062 579134
rect 578146 578898 578382 579134
rect 577826 543218 578062 543454
rect 578146 543218 578382 543454
rect 577826 542898 578062 543134
rect 578146 542898 578382 543134
rect 577826 507218 578062 507454
rect 578146 507218 578382 507454
rect 577826 506898 578062 507134
rect 578146 506898 578382 507134
rect 577826 471218 578062 471454
rect 578146 471218 578382 471454
rect 577826 470898 578062 471134
rect 578146 470898 578382 471134
rect 577826 435218 578062 435454
rect 578146 435218 578382 435454
rect 577826 434898 578062 435134
rect 578146 434898 578382 435134
rect 577826 399218 578062 399454
rect 578146 399218 578382 399454
rect 577826 398898 578062 399134
rect 578146 398898 578382 399134
rect 577826 363218 578062 363454
rect 578146 363218 578382 363454
rect 577826 362898 578062 363134
rect 578146 362898 578382 363134
rect 577826 327218 578062 327454
rect 578146 327218 578382 327454
rect 577826 326898 578062 327134
rect 578146 326898 578382 327134
rect 577826 291218 578062 291454
rect 578146 291218 578382 291454
rect 577826 290898 578062 291134
rect 578146 290898 578382 291134
rect 577826 255218 578062 255454
rect 578146 255218 578382 255454
rect 577826 254898 578062 255134
rect 578146 254898 578382 255134
rect 577826 219218 578062 219454
rect 578146 219218 578382 219454
rect 577826 218898 578062 219134
rect 578146 218898 578382 219134
rect 577826 183218 578062 183454
rect 578146 183218 578382 183454
rect 577826 182898 578062 183134
rect 578146 182898 578382 183134
rect 577826 147218 578062 147454
rect 578146 147218 578382 147454
rect 577826 146898 578062 147134
rect 578146 146898 578382 147134
rect 577826 111218 578062 111454
rect 578146 111218 578382 111454
rect 577826 110898 578062 111134
rect 578146 110898 578382 111134
rect 577826 75218 578062 75454
rect 578146 75218 578382 75454
rect 577826 74898 578062 75134
rect 578146 74898 578382 75134
rect 577826 39218 578062 39454
rect 578146 39218 578382 39454
rect 577826 38898 578062 39134
rect 578146 38898 578382 39134
rect 577826 3218 578062 3454
rect 578146 3218 578382 3454
rect 577826 2898 578062 3134
rect 578146 2898 578382 3134
rect 577826 -582 578062 -346
rect 578146 -582 578382 -346
rect 577826 -902 578062 -666
rect 578146 -902 578382 -666
rect 587262 706522 587498 706758
rect 587582 706522 587818 706758
rect 587262 706202 587498 706438
rect 587582 706202 587818 706438
rect 586302 705562 586538 705798
rect 586622 705562 586858 705798
rect 586302 705242 586538 705478
rect 586622 705242 586858 705478
rect 581546 690938 581782 691174
rect 581866 690938 582102 691174
rect 581546 690618 581782 690854
rect 581866 690618 582102 690854
rect 581546 654938 581782 655174
rect 581866 654938 582102 655174
rect 581546 654618 581782 654854
rect 581866 654618 582102 654854
rect 581546 618938 581782 619174
rect 581866 618938 582102 619174
rect 581546 618618 581782 618854
rect 581866 618618 582102 618854
rect 581546 582938 581782 583174
rect 581866 582938 582102 583174
rect 581546 582618 581782 582854
rect 581866 582618 582102 582854
rect 581546 546938 581782 547174
rect 581866 546938 582102 547174
rect 581546 546618 581782 546854
rect 581866 546618 582102 546854
rect 581546 510938 581782 511174
rect 581866 510938 582102 511174
rect 581546 510618 581782 510854
rect 581866 510618 582102 510854
rect 581546 474938 581782 475174
rect 581866 474938 582102 475174
rect 581546 474618 581782 474854
rect 581866 474618 582102 474854
rect 581546 438938 581782 439174
rect 581866 438938 582102 439174
rect 581546 438618 581782 438854
rect 581866 438618 582102 438854
rect 581546 402938 581782 403174
rect 581866 402938 582102 403174
rect 581546 402618 581782 402854
rect 581866 402618 582102 402854
rect 581546 366938 581782 367174
rect 581866 366938 582102 367174
rect 581546 366618 581782 366854
rect 581866 366618 582102 366854
rect 581546 330938 581782 331174
rect 581866 330938 582102 331174
rect 581546 330618 581782 330854
rect 581866 330618 582102 330854
rect 581546 294938 581782 295174
rect 581866 294938 582102 295174
rect 581546 294618 581782 294854
rect 581866 294618 582102 294854
rect 581546 258938 581782 259174
rect 581866 258938 582102 259174
rect 581546 258618 581782 258854
rect 581866 258618 582102 258854
rect 581546 222938 581782 223174
rect 581866 222938 582102 223174
rect 581546 222618 581782 222854
rect 581866 222618 582102 222854
rect 581546 186938 581782 187174
rect 581866 186938 582102 187174
rect 581546 186618 581782 186854
rect 581866 186618 582102 186854
rect 581546 150938 581782 151174
rect 581866 150938 582102 151174
rect 581546 150618 581782 150854
rect 581866 150618 582102 150854
rect 581546 114938 581782 115174
rect 581866 114938 582102 115174
rect 581546 114618 581782 114854
rect 581866 114618 582102 114854
rect 581546 78938 581782 79174
rect 581866 78938 582102 79174
rect 581546 78618 581782 78854
rect 581866 78618 582102 78854
rect 581546 42938 581782 43174
rect 581866 42938 582102 43174
rect 581546 42618 581782 42854
rect 581866 42618 582102 42854
rect 581546 6938 581782 7174
rect 581866 6938 582102 7174
rect 581546 6618 581782 6854
rect 581866 6618 582102 6854
rect 585342 704602 585578 704838
rect 585662 704602 585898 704838
rect 585342 704282 585578 704518
rect 585662 704282 585898 704518
rect 585342 687218 585578 687454
rect 585662 687218 585898 687454
rect 585342 686898 585578 687134
rect 585662 686898 585898 687134
rect 585342 651218 585578 651454
rect 585662 651218 585898 651454
rect 585342 650898 585578 651134
rect 585662 650898 585898 651134
rect 585342 615218 585578 615454
rect 585662 615218 585898 615454
rect 585342 614898 585578 615134
rect 585662 614898 585898 615134
rect 585342 579218 585578 579454
rect 585662 579218 585898 579454
rect 585342 578898 585578 579134
rect 585662 578898 585898 579134
rect 585342 543218 585578 543454
rect 585662 543218 585898 543454
rect 585342 542898 585578 543134
rect 585662 542898 585898 543134
rect 585342 507218 585578 507454
rect 585662 507218 585898 507454
rect 585342 506898 585578 507134
rect 585662 506898 585898 507134
rect 585342 471218 585578 471454
rect 585662 471218 585898 471454
rect 585342 470898 585578 471134
rect 585662 470898 585898 471134
rect 585342 435218 585578 435454
rect 585662 435218 585898 435454
rect 585342 434898 585578 435134
rect 585662 434898 585898 435134
rect 585342 399218 585578 399454
rect 585662 399218 585898 399454
rect 585342 398898 585578 399134
rect 585662 398898 585898 399134
rect 585342 363218 585578 363454
rect 585662 363218 585898 363454
rect 585342 362898 585578 363134
rect 585662 362898 585898 363134
rect 585342 327218 585578 327454
rect 585662 327218 585898 327454
rect 585342 326898 585578 327134
rect 585662 326898 585898 327134
rect 585342 291218 585578 291454
rect 585662 291218 585898 291454
rect 585342 290898 585578 291134
rect 585662 290898 585898 291134
rect 585342 255218 585578 255454
rect 585662 255218 585898 255454
rect 585342 254898 585578 255134
rect 585662 254898 585898 255134
rect 585342 219218 585578 219454
rect 585662 219218 585898 219454
rect 585342 218898 585578 219134
rect 585662 218898 585898 219134
rect 585342 183218 585578 183454
rect 585662 183218 585898 183454
rect 585342 182898 585578 183134
rect 585662 182898 585898 183134
rect 585342 147218 585578 147454
rect 585662 147218 585898 147454
rect 585342 146898 585578 147134
rect 585662 146898 585898 147134
rect 585342 111218 585578 111454
rect 585662 111218 585898 111454
rect 585342 110898 585578 111134
rect 585662 110898 585898 111134
rect 585342 75218 585578 75454
rect 585662 75218 585898 75454
rect 585342 74898 585578 75134
rect 585662 74898 585898 75134
rect 585342 39218 585578 39454
rect 585662 39218 585898 39454
rect 585342 38898 585578 39134
rect 585662 38898 585898 39134
rect 585342 3218 585578 3454
rect 585662 3218 585898 3454
rect 585342 2898 585578 3134
rect 585662 2898 585898 3134
rect 585342 -582 585578 -346
rect 585662 -582 585898 -346
rect 585342 -902 585578 -666
rect 585662 -902 585898 -666
rect 586302 669218 586538 669454
rect 586622 669218 586858 669454
rect 586302 668898 586538 669134
rect 586622 668898 586858 669134
rect 586302 633218 586538 633454
rect 586622 633218 586858 633454
rect 586302 632898 586538 633134
rect 586622 632898 586858 633134
rect 586302 597218 586538 597454
rect 586622 597218 586858 597454
rect 586302 596898 586538 597134
rect 586622 596898 586858 597134
rect 586302 561218 586538 561454
rect 586622 561218 586858 561454
rect 586302 560898 586538 561134
rect 586622 560898 586858 561134
rect 586302 525218 586538 525454
rect 586622 525218 586858 525454
rect 586302 524898 586538 525134
rect 586622 524898 586858 525134
rect 586302 489218 586538 489454
rect 586622 489218 586858 489454
rect 586302 488898 586538 489134
rect 586622 488898 586858 489134
rect 586302 453218 586538 453454
rect 586622 453218 586858 453454
rect 586302 452898 586538 453134
rect 586622 452898 586858 453134
rect 586302 417218 586538 417454
rect 586622 417218 586858 417454
rect 586302 416898 586538 417134
rect 586622 416898 586858 417134
rect 586302 381218 586538 381454
rect 586622 381218 586858 381454
rect 586302 380898 586538 381134
rect 586622 380898 586858 381134
rect 586302 345218 586538 345454
rect 586622 345218 586858 345454
rect 586302 344898 586538 345134
rect 586622 344898 586858 345134
rect 586302 309218 586538 309454
rect 586622 309218 586858 309454
rect 586302 308898 586538 309134
rect 586622 308898 586858 309134
rect 586302 273218 586538 273454
rect 586622 273218 586858 273454
rect 586302 272898 586538 273134
rect 586622 272898 586858 273134
rect 586302 237218 586538 237454
rect 586622 237218 586858 237454
rect 586302 236898 586538 237134
rect 586622 236898 586858 237134
rect 586302 201218 586538 201454
rect 586622 201218 586858 201454
rect 586302 200898 586538 201134
rect 586622 200898 586858 201134
rect 586302 165218 586538 165454
rect 586622 165218 586858 165454
rect 586302 164898 586538 165134
rect 586622 164898 586858 165134
rect 586302 129218 586538 129454
rect 586622 129218 586858 129454
rect 586302 128898 586538 129134
rect 586622 128898 586858 129134
rect 586302 93218 586538 93454
rect 586622 93218 586858 93454
rect 586302 92898 586538 93134
rect 586622 92898 586858 93134
rect 586302 57218 586538 57454
rect 586622 57218 586858 57454
rect 586302 56898 586538 57134
rect 586622 56898 586858 57134
rect 586302 21218 586538 21454
rect 586622 21218 586858 21454
rect 586302 20898 586538 21134
rect 586622 20898 586858 21134
rect 586302 -1542 586538 -1306
rect 586622 -1542 586858 -1306
rect 586302 -1862 586538 -1626
rect 586622 -1862 586858 -1626
rect 587262 690938 587498 691174
rect 587582 690938 587818 691174
rect 587262 690618 587498 690854
rect 587582 690618 587818 690854
rect 587262 654938 587498 655174
rect 587582 654938 587818 655174
rect 587262 654618 587498 654854
rect 587582 654618 587818 654854
rect 587262 618938 587498 619174
rect 587582 618938 587818 619174
rect 587262 618618 587498 618854
rect 587582 618618 587818 618854
rect 587262 582938 587498 583174
rect 587582 582938 587818 583174
rect 587262 582618 587498 582854
rect 587582 582618 587818 582854
rect 587262 546938 587498 547174
rect 587582 546938 587818 547174
rect 587262 546618 587498 546854
rect 587582 546618 587818 546854
rect 587262 510938 587498 511174
rect 587582 510938 587818 511174
rect 587262 510618 587498 510854
rect 587582 510618 587818 510854
rect 587262 474938 587498 475174
rect 587582 474938 587818 475174
rect 587262 474618 587498 474854
rect 587582 474618 587818 474854
rect 587262 438938 587498 439174
rect 587582 438938 587818 439174
rect 587262 438618 587498 438854
rect 587582 438618 587818 438854
rect 587262 402938 587498 403174
rect 587582 402938 587818 403174
rect 587262 402618 587498 402854
rect 587582 402618 587818 402854
rect 587262 366938 587498 367174
rect 587582 366938 587818 367174
rect 587262 366618 587498 366854
rect 587582 366618 587818 366854
rect 587262 330938 587498 331174
rect 587582 330938 587818 331174
rect 587262 330618 587498 330854
rect 587582 330618 587818 330854
rect 587262 294938 587498 295174
rect 587582 294938 587818 295174
rect 587262 294618 587498 294854
rect 587582 294618 587818 294854
rect 587262 258938 587498 259174
rect 587582 258938 587818 259174
rect 587262 258618 587498 258854
rect 587582 258618 587818 258854
rect 587262 222938 587498 223174
rect 587582 222938 587818 223174
rect 587262 222618 587498 222854
rect 587582 222618 587818 222854
rect 587262 186938 587498 187174
rect 587582 186938 587818 187174
rect 587262 186618 587498 186854
rect 587582 186618 587818 186854
rect 587262 150938 587498 151174
rect 587582 150938 587818 151174
rect 587262 150618 587498 150854
rect 587582 150618 587818 150854
rect 587262 114938 587498 115174
rect 587582 114938 587818 115174
rect 587262 114618 587498 114854
rect 587582 114618 587818 114854
rect 587262 78938 587498 79174
rect 587582 78938 587818 79174
rect 587262 78618 587498 78854
rect 587582 78618 587818 78854
rect 587262 42938 587498 43174
rect 587582 42938 587818 43174
rect 587262 42618 587498 42854
rect 587582 42618 587818 42854
rect 587262 6938 587498 7174
rect 587582 6938 587818 7174
rect 587262 6618 587498 6854
rect 587582 6618 587818 6854
rect 581546 -2502 581782 -2266
rect 581866 -2502 582102 -2266
rect 581546 -2822 581782 -2586
rect 581866 -2822 582102 -2586
rect 587262 -2502 587498 -2266
rect 587582 -2502 587818 -2266
rect 587262 -2822 587498 -2586
rect 587582 -2822 587818 -2586
rect 588222 672938 588458 673174
rect 588542 672938 588778 673174
rect 588222 672618 588458 672854
rect 588542 672618 588778 672854
rect 588222 636938 588458 637174
rect 588542 636938 588778 637174
rect 588222 636618 588458 636854
rect 588542 636618 588778 636854
rect 588222 600938 588458 601174
rect 588542 600938 588778 601174
rect 588222 600618 588458 600854
rect 588542 600618 588778 600854
rect 588222 564938 588458 565174
rect 588542 564938 588778 565174
rect 588222 564618 588458 564854
rect 588542 564618 588778 564854
rect 588222 528938 588458 529174
rect 588542 528938 588778 529174
rect 588222 528618 588458 528854
rect 588542 528618 588778 528854
rect 588222 492938 588458 493174
rect 588542 492938 588778 493174
rect 588222 492618 588458 492854
rect 588542 492618 588778 492854
rect 588222 456938 588458 457174
rect 588542 456938 588778 457174
rect 588222 456618 588458 456854
rect 588542 456618 588778 456854
rect 588222 420938 588458 421174
rect 588542 420938 588778 421174
rect 588222 420618 588458 420854
rect 588542 420618 588778 420854
rect 588222 384938 588458 385174
rect 588542 384938 588778 385174
rect 588222 384618 588458 384854
rect 588542 384618 588778 384854
rect 588222 348938 588458 349174
rect 588542 348938 588778 349174
rect 588222 348618 588458 348854
rect 588542 348618 588778 348854
rect 588222 312938 588458 313174
rect 588542 312938 588778 313174
rect 588222 312618 588458 312854
rect 588542 312618 588778 312854
rect 588222 276938 588458 277174
rect 588542 276938 588778 277174
rect 588222 276618 588458 276854
rect 588542 276618 588778 276854
rect 588222 240938 588458 241174
rect 588542 240938 588778 241174
rect 588222 240618 588458 240854
rect 588542 240618 588778 240854
rect 588222 204938 588458 205174
rect 588542 204938 588778 205174
rect 588222 204618 588458 204854
rect 588542 204618 588778 204854
rect 588222 168938 588458 169174
rect 588542 168938 588778 169174
rect 588222 168618 588458 168854
rect 588542 168618 588778 168854
rect 588222 132938 588458 133174
rect 588542 132938 588778 133174
rect 588222 132618 588458 132854
rect 588542 132618 588778 132854
rect 588222 96938 588458 97174
rect 588542 96938 588778 97174
rect 588222 96618 588458 96854
rect 588542 96618 588778 96854
rect 588222 60938 588458 61174
rect 588542 60938 588778 61174
rect 588222 60618 588458 60854
rect 588542 60618 588778 60854
rect 588222 24938 588458 25174
rect 588542 24938 588778 25174
rect 588222 24618 588458 24854
rect 588542 24618 588778 24854
rect 588222 -3462 588458 -3226
rect 588542 -3462 588778 -3226
rect 588222 -3782 588458 -3546
rect 588542 -3782 588778 -3546
rect 589182 694658 589418 694894
rect 589502 694658 589738 694894
rect 589182 694338 589418 694574
rect 589502 694338 589738 694574
rect 589182 658658 589418 658894
rect 589502 658658 589738 658894
rect 589182 658338 589418 658574
rect 589502 658338 589738 658574
rect 589182 622658 589418 622894
rect 589502 622658 589738 622894
rect 589182 622338 589418 622574
rect 589502 622338 589738 622574
rect 589182 586658 589418 586894
rect 589502 586658 589738 586894
rect 589182 586338 589418 586574
rect 589502 586338 589738 586574
rect 589182 550658 589418 550894
rect 589502 550658 589738 550894
rect 589182 550338 589418 550574
rect 589502 550338 589738 550574
rect 589182 514658 589418 514894
rect 589502 514658 589738 514894
rect 589182 514338 589418 514574
rect 589502 514338 589738 514574
rect 589182 478658 589418 478894
rect 589502 478658 589738 478894
rect 589182 478338 589418 478574
rect 589502 478338 589738 478574
rect 589182 442658 589418 442894
rect 589502 442658 589738 442894
rect 589182 442338 589418 442574
rect 589502 442338 589738 442574
rect 589182 406658 589418 406894
rect 589502 406658 589738 406894
rect 589182 406338 589418 406574
rect 589502 406338 589738 406574
rect 589182 370658 589418 370894
rect 589502 370658 589738 370894
rect 589182 370338 589418 370574
rect 589502 370338 589738 370574
rect 589182 334658 589418 334894
rect 589502 334658 589738 334894
rect 589182 334338 589418 334574
rect 589502 334338 589738 334574
rect 589182 298658 589418 298894
rect 589502 298658 589738 298894
rect 589182 298338 589418 298574
rect 589502 298338 589738 298574
rect 589182 262658 589418 262894
rect 589502 262658 589738 262894
rect 589182 262338 589418 262574
rect 589502 262338 589738 262574
rect 589182 226658 589418 226894
rect 589502 226658 589738 226894
rect 589182 226338 589418 226574
rect 589502 226338 589738 226574
rect 589182 190658 589418 190894
rect 589502 190658 589738 190894
rect 589182 190338 589418 190574
rect 589502 190338 589738 190574
rect 589182 154658 589418 154894
rect 589502 154658 589738 154894
rect 589182 154338 589418 154574
rect 589502 154338 589738 154574
rect 589182 118658 589418 118894
rect 589502 118658 589738 118894
rect 589182 118338 589418 118574
rect 589502 118338 589738 118574
rect 589182 82658 589418 82894
rect 589502 82658 589738 82894
rect 589182 82338 589418 82574
rect 589502 82338 589738 82574
rect 589182 46658 589418 46894
rect 589502 46658 589738 46894
rect 589182 46338 589418 46574
rect 589502 46338 589738 46574
rect 589182 10658 589418 10894
rect 589502 10658 589738 10894
rect 589182 10338 589418 10574
rect 589502 10338 589738 10574
rect 589182 -4422 589418 -4186
rect 589502 -4422 589738 -4186
rect 589182 -4742 589418 -4506
rect 589502 -4742 589738 -4506
rect 590142 676658 590378 676894
rect 590462 676658 590698 676894
rect 590142 676338 590378 676574
rect 590462 676338 590698 676574
rect 590142 640658 590378 640894
rect 590462 640658 590698 640894
rect 590142 640338 590378 640574
rect 590462 640338 590698 640574
rect 590142 604658 590378 604894
rect 590462 604658 590698 604894
rect 590142 604338 590378 604574
rect 590462 604338 590698 604574
rect 590142 568658 590378 568894
rect 590462 568658 590698 568894
rect 590142 568338 590378 568574
rect 590462 568338 590698 568574
rect 590142 532658 590378 532894
rect 590462 532658 590698 532894
rect 590142 532338 590378 532574
rect 590462 532338 590698 532574
rect 590142 496658 590378 496894
rect 590462 496658 590698 496894
rect 590142 496338 590378 496574
rect 590462 496338 590698 496574
rect 590142 460658 590378 460894
rect 590462 460658 590698 460894
rect 590142 460338 590378 460574
rect 590462 460338 590698 460574
rect 590142 424658 590378 424894
rect 590462 424658 590698 424894
rect 590142 424338 590378 424574
rect 590462 424338 590698 424574
rect 590142 388658 590378 388894
rect 590462 388658 590698 388894
rect 590142 388338 590378 388574
rect 590462 388338 590698 388574
rect 590142 352658 590378 352894
rect 590462 352658 590698 352894
rect 590142 352338 590378 352574
rect 590462 352338 590698 352574
rect 590142 316658 590378 316894
rect 590462 316658 590698 316894
rect 590142 316338 590378 316574
rect 590462 316338 590698 316574
rect 590142 280658 590378 280894
rect 590462 280658 590698 280894
rect 590142 280338 590378 280574
rect 590462 280338 590698 280574
rect 590142 244658 590378 244894
rect 590462 244658 590698 244894
rect 590142 244338 590378 244574
rect 590462 244338 590698 244574
rect 590142 208658 590378 208894
rect 590462 208658 590698 208894
rect 590142 208338 590378 208574
rect 590462 208338 590698 208574
rect 590142 172658 590378 172894
rect 590462 172658 590698 172894
rect 590142 172338 590378 172574
rect 590462 172338 590698 172574
rect 590142 136658 590378 136894
rect 590462 136658 590698 136894
rect 590142 136338 590378 136574
rect 590462 136338 590698 136574
rect 590142 100658 590378 100894
rect 590462 100658 590698 100894
rect 590142 100338 590378 100574
rect 590462 100338 590698 100574
rect 590142 64658 590378 64894
rect 590462 64658 590698 64894
rect 590142 64338 590378 64574
rect 590462 64338 590698 64574
rect 590142 28658 590378 28894
rect 590462 28658 590698 28894
rect 590142 28338 590378 28574
rect 590462 28338 590698 28574
rect 590142 -5382 590378 -5146
rect 590462 -5382 590698 -5146
rect 590142 -5702 590378 -5466
rect 590462 -5702 590698 -5466
rect 591102 698378 591338 698614
rect 591422 698378 591658 698614
rect 591102 698058 591338 698294
rect 591422 698058 591658 698294
rect 591102 662378 591338 662614
rect 591422 662378 591658 662614
rect 591102 662058 591338 662294
rect 591422 662058 591658 662294
rect 591102 626378 591338 626614
rect 591422 626378 591658 626614
rect 591102 626058 591338 626294
rect 591422 626058 591658 626294
rect 591102 590378 591338 590614
rect 591422 590378 591658 590614
rect 591102 590058 591338 590294
rect 591422 590058 591658 590294
rect 591102 554378 591338 554614
rect 591422 554378 591658 554614
rect 591102 554058 591338 554294
rect 591422 554058 591658 554294
rect 591102 518378 591338 518614
rect 591422 518378 591658 518614
rect 591102 518058 591338 518294
rect 591422 518058 591658 518294
rect 591102 482378 591338 482614
rect 591422 482378 591658 482614
rect 591102 482058 591338 482294
rect 591422 482058 591658 482294
rect 591102 446378 591338 446614
rect 591422 446378 591658 446614
rect 591102 446058 591338 446294
rect 591422 446058 591658 446294
rect 591102 410378 591338 410614
rect 591422 410378 591658 410614
rect 591102 410058 591338 410294
rect 591422 410058 591658 410294
rect 591102 374378 591338 374614
rect 591422 374378 591658 374614
rect 591102 374058 591338 374294
rect 591422 374058 591658 374294
rect 591102 338378 591338 338614
rect 591422 338378 591658 338614
rect 591102 338058 591338 338294
rect 591422 338058 591658 338294
rect 591102 302378 591338 302614
rect 591422 302378 591658 302614
rect 591102 302058 591338 302294
rect 591422 302058 591658 302294
rect 591102 266378 591338 266614
rect 591422 266378 591658 266614
rect 591102 266058 591338 266294
rect 591422 266058 591658 266294
rect 591102 230378 591338 230614
rect 591422 230378 591658 230614
rect 591102 230058 591338 230294
rect 591422 230058 591658 230294
rect 591102 194378 591338 194614
rect 591422 194378 591658 194614
rect 591102 194058 591338 194294
rect 591422 194058 591658 194294
rect 591102 158378 591338 158614
rect 591422 158378 591658 158614
rect 591102 158058 591338 158294
rect 591422 158058 591658 158294
rect 591102 122378 591338 122614
rect 591422 122378 591658 122614
rect 591102 122058 591338 122294
rect 591422 122058 591658 122294
rect 591102 86378 591338 86614
rect 591422 86378 591658 86614
rect 591102 86058 591338 86294
rect 591422 86058 591658 86294
rect 591102 50378 591338 50614
rect 591422 50378 591658 50614
rect 591102 50058 591338 50294
rect 591422 50058 591658 50294
rect 591102 14378 591338 14614
rect 591422 14378 591658 14614
rect 591102 14058 591338 14294
rect 591422 14058 591658 14294
rect 591102 -6342 591338 -6106
rect 591422 -6342 591658 -6106
rect 591102 -6662 591338 -6426
rect 591422 -6662 591658 -6426
rect 592062 680378 592298 680614
rect 592382 680378 592618 680614
rect 592062 680058 592298 680294
rect 592382 680058 592618 680294
rect 592062 644378 592298 644614
rect 592382 644378 592618 644614
rect 592062 644058 592298 644294
rect 592382 644058 592618 644294
rect 592062 608378 592298 608614
rect 592382 608378 592618 608614
rect 592062 608058 592298 608294
rect 592382 608058 592618 608294
rect 592062 572378 592298 572614
rect 592382 572378 592618 572614
rect 592062 572058 592298 572294
rect 592382 572058 592618 572294
rect 592062 536378 592298 536614
rect 592382 536378 592618 536614
rect 592062 536058 592298 536294
rect 592382 536058 592618 536294
rect 592062 500378 592298 500614
rect 592382 500378 592618 500614
rect 592062 500058 592298 500294
rect 592382 500058 592618 500294
rect 592062 464378 592298 464614
rect 592382 464378 592618 464614
rect 592062 464058 592298 464294
rect 592382 464058 592618 464294
rect 592062 428378 592298 428614
rect 592382 428378 592618 428614
rect 592062 428058 592298 428294
rect 592382 428058 592618 428294
rect 592062 392378 592298 392614
rect 592382 392378 592618 392614
rect 592062 392058 592298 392294
rect 592382 392058 592618 392294
rect 592062 356378 592298 356614
rect 592382 356378 592618 356614
rect 592062 356058 592298 356294
rect 592382 356058 592618 356294
rect 592062 320378 592298 320614
rect 592382 320378 592618 320614
rect 592062 320058 592298 320294
rect 592382 320058 592618 320294
rect 592062 284378 592298 284614
rect 592382 284378 592618 284614
rect 592062 284058 592298 284294
rect 592382 284058 592618 284294
rect 592062 248378 592298 248614
rect 592382 248378 592618 248614
rect 592062 248058 592298 248294
rect 592382 248058 592618 248294
rect 592062 212378 592298 212614
rect 592382 212378 592618 212614
rect 592062 212058 592298 212294
rect 592382 212058 592618 212294
rect 592062 176378 592298 176614
rect 592382 176378 592618 176614
rect 592062 176058 592298 176294
rect 592382 176058 592618 176294
rect 592062 140378 592298 140614
rect 592382 140378 592618 140614
rect 592062 140058 592298 140294
rect 592382 140058 592618 140294
rect 592062 104378 592298 104614
rect 592382 104378 592618 104614
rect 592062 104058 592298 104294
rect 592382 104058 592618 104294
rect 592062 68378 592298 68614
rect 592382 68378 592618 68614
rect 592062 68058 592298 68294
rect 592382 68058 592618 68294
rect 592062 32378 592298 32614
rect 592382 32378 592618 32614
rect 592062 32058 592298 32294
rect 592382 32058 592618 32294
rect 570986 -7302 571222 -7066
rect 571306 -7302 571542 -7066
rect 570986 -7622 571222 -7386
rect 571306 -7622 571542 -7386
rect 592062 -7302 592298 -7066
rect 592382 -7302 592618 -7066
rect 592062 -7622 592298 -7386
rect 592382 -7622 592618 -7386
<< metal5 >>
rect -8726 711558 592650 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 30986 711558
rect 31222 711322 31306 711558
rect 31542 711322 66986 711558
rect 67222 711322 67306 711558
rect 67542 711322 102986 711558
rect 103222 711322 103306 711558
rect 103542 711322 138986 711558
rect 139222 711322 139306 711558
rect 139542 711322 174986 711558
rect 175222 711322 175306 711558
rect 175542 711322 210986 711558
rect 211222 711322 211306 711558
rect 211542 711322 246986 711558
rect 247222 711322 247306 711558
rect 247542 711322 282986 711558
rect 283222 711322 283306 711558
rect 283542 711322 318986 711558
rect 319222 711322 319306 711558
rect 319542 711322 354986 711558
rect 355222 711322 355306 711558
rect 355542 711322 390986 711558
rect 391222 711322 391306 711558
rect 391542 711322 426986 711558
rect 427222 711322 427306 711558
rect 427542 711322 462986 711558
rect 463222 711322 463306 711558
rect 463542 711322 498986 711558
rect 499222 711322 499306 711558
rect 499542 711322 534986 711558
rect 535222 711322 535306 711558
rect 535542 711322 570986 711558
rect 571222 711322 571306 711558
rect 571542 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect -8726 711238 592650 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 30986 711238
rect 31222 711002 31306 711238
rect 31542 711002 66986 711238
rect 67222 711002 67306 711238
rect 67542 711002 102986 711238
rect 103222 711002 103306 711238
rect 103542 711002 138986 711238
rect 139222 711002 139306 711238
rect 139542 711002 174986 711238
rect 175222 711002 175306 711238
rect 175542 711002 210986 711238
rect 211222 711002 211306 711238
rect 211542 711002 246986 711238
rect 247222 711002 247306 711238
rect 247542 711002 282986 711238
rect 283222 711002 283306 711238
rect 283542 711002 318986 711238
rect 319222 711002 319306 711238
rect 319542 711002 354986 711238
rect 355222 711002 355306 711238
rect 355542 711002 390986 711238
rect 391222 711002 391306 711238
rect 391542 711002 426986 711238
rect 427222 711002 427306 711238
rect 427542 711002 462986 711238
rect 463222 711002 463306 711238
rect 463542 711002 498986 711238
rect 499222 711002 499306 711238
rect 499542 711002 534986 711238
rect 535222 711002 535306 711238
rect 535542 711002 570986 711238
rect 571222 711002 571306 711238
rect 571542 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect -8726 710970 592650 711002
rect -7766 710598 591690 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 12986 710598
rect 13222 710362 13306 710598
rect 13542 710362 48986 710598
rect 49222 710362 49306 710598
rect 49542 710362 84986 710598
rect 85222 710362 85306 710598
rect 85542 710362 120986 710598
rect 121222 710362 121306 710598
rect 121542 710362 156986 710598
rect 157222 710362 157306 710598
rect 157542 710362 192986 710598
rect 193222 710362 193306 710598
rect 193542 710362 228986 710598
rect 229222 710362 229306 710598
rect 229542 710362 264986 710598
rect 265222 710362 265306 710598
rect 265542 710362 300986 710598
rect 301222 710362 301306 710598
rect 301542 710362 336986 710598
rect 337222 710362 337306 710598
rect 337542 710362 372986 710598
rect 373222 710362 373306 710598
rect 373542 710362 408986 710598
rect 409222 710362 409306 710598
rect 409542 710362 444986 710598
rect 445222 710362 445306 710598
rect 445542 710362 480986 710598
rect 481222 710362 481306 710598
rect 481542 710362 516986 710598
rect 517222 710362 517306 710598
rect 517542 710362 552986 710598
rect 553222 710362 553306 710598
rect 553542 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect -7766 710278 591690 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 12986 710278
rect 13222 710042 13306 710278
rect 13542 710042 48986 710278
rect 49222 710042 49306 710278
rect 49542 710042 84986 710278
rect 85222 710042 85306 710278
rect 85542 710042 120986 710278
rect 121222 710042 121306 710278
rect 121542 710042 156986 710278
rect 157222 710042 157306 710278
rect 157542 710042 192986 710278
rect 193222 710042 193306 710278
rect 193542 710042 228986 710278
rect 229222 710042 229306 710278
rect 229542 710042 264986 710278
rect 265222 710042 265306 710278
rect 265542 710042 300986 710278
rect 301222 710042 301306 710278
rect 301542 710042 336986 710278
rect 337222 710042 337306 710278
rect 337542 710042 372986 710278
rect 373222 710042 373306 710278
rect 373542 710042 408986 710278
rect 409222 710042 409306 710278
rect 409542 710042 444986 710278
rect 445222 710042 445306 710278
rect 445542 710042 480986 710278
rect 481222 710042 481306 710278
rect 481542 710042 516986 710278
rect 517222 710042 517306 710278
rect 517542 710042 552986 710278
rect 553222 710042 553306 710278
rect 553542 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect -7766 710010 591690 710042
rect -6806 709638 590730 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 27266 709638
rect 27502 709402 27586 709638
rect 27822 709402 63266 709638
rect 63502 709402 63586 709638
rect 63822 709402 99266 709638
rect 99502 709402 99586 709638
rect 99822 709402 135266 709638
rect 135502 709402 135586 709638
rect 135822 709402 171266 709638
rect 171502 709402 171586 709638
rect 171822 709402 207266 709638
rect 207502 709402 207586 709638
rect 207822 709402 243266 709638
rect 243502 709402 243586 709638
rect 243822 709402 279266 709638
rect 279502 709402 279586 709638
rect 279822 709402 315266 709638
rect 315502 709402 315586 709638
rect 315822 709402 351266 709638
rect 351502 709402 351586 709638
rect 351822 709402 387266 709638
rect 387502 709402 387586 709638
rect 387822 709402 423266 709638
rect 423502 709402 423586 709638
rect 423822 709402 459266 709638
rect 459502 709402 459586 709638
rect 459822 709402 495266 709638
rect 495502 709402 495586 709638
rect 495822 709402 531266 709638
rect 531502 709402 531586 709638
rect 531822 709402 567266 709638
rect 567502 709402 567586 709638
rect 567822 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect -6806 709318 590730 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 27266 709318
rect 27502 709082 27586 709318
rect 27822 709082 63266 709318
rect 63502 709082 63586 709318
rect 63822 709082 99266 709318
rect 99502 709082 99586 709318
rect 99822 709082 135266 709318
rect 135502 709082 135586 709318
rect 135822 709082 171266 709318
rect 171502 709082 171586 709318
rect 171822 709082 207266 709318
rect 207502 709082 207586 709318
rect 207822 709082 243266 709318
rect 243502 709082 243586 709318
rect 243822 709082 279266 709318
rect 279502 709082 279586 709318
rect 279822 709082 315266 709318
rect 315502 709082 315586 709318
rect 315822 709082 351266 709318
rect 351502 709082 351586 709318
rect 351822 709082 387266 709318
rect 387502 709082 387586 709318
rect 387822 709082 423266 709318
rect 423502 709082 423586 709318
rect 423822 709082 459266 709318
rect 459502 709082 459586 709318
rect 459822 709082 495266 709318
rect 495502 709082 495586 709318
rect 495822 709082 531266 709318
rect 531502 709082 531586 709318
rect 531822 709082 567266 709318
rect 567502 709082 567586 709318
rect 567822 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect -6806 709050 590730 709082
rect -5846 708678 589770 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 9266 708678
rect 9502 708442 9586 708678
rect 9822 708442 45266 708678
rect 45502 708442 45586 708678
rect 45822 708442 81266 708678
rect 81502 708442 81586 708678
rect 81822 708442 117266 708678
rect 117502 708442 117586 708678
rect 117822 708442 153266 708678
rect 153502 708442 153586 708678
rect 153822 708442 189266 708678
rect 189502 708442 189586 708678
rect 189822 708442 225266 708678
rect 225502 708442 225586 708678
rect 225822 708442 261266 708678
rect 261502 708442 261586 708678
rect 261822 708442 297266 708678
rect 297502 708442 297586 708678
rect 297822 708442 333266 708678
rect 333502 708442 333586 708678
rect 333822 708442 369266 708678
rect 369502 708442 369586 708678
rect 369822 708442 405266 708678
rect 405502 708442 405586 708678
rect 405822 708442 441266 708678
rect 441502 708442 441586 708678
rect 441822 708442 477266 708678
rect 477502 708442 477586 708678
rect 477822 708442 513266 708678
rect 513502 708442 513586 708678
rect 513822 708442 549266 708678
rect 549502 708442 549586 708678
rect 549822 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect -5846 708358 589770 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 9266 708358
rect 9502 708122 9586 708358
rect 9822 708122 45266 708358
rect 45502 708122 45586 708358
rect 45822 708122 81266 708358
rect 81502 708122 81586 708358
rect 81822 708122 117266 708358
rect 117502 708122 117586 708358
rect 117822 708122 153266 708358
rect 153502 708122 153586 708358
rect 153822 708122 189266 708358
rect 189502 708122 189586 708358
rect 189822 708122 225266 708358
rect 225502 708122 225586 708358
rect 225822 708122 261266 708358
rect 261502 708122 261586 708358
rect 261822 708122 297266 708358
rect 297502 708122 297586 708358
rect 297822 708122 333266 708358
rect 333502 708122 333586 708358
rect 333822 708122 369266 708358
rect 369502 708122 369586 708358
rect 369822 708122 405266 708358
rect 405502 708122 405586 708358
rect 405822 708122 441266 708358
rect 441502 708122 441586 708358
rect 441822 708122 477266 708358
rect 477502 708122 477586 708358
rect 477822 708122 513266 708358
rect 513502 708122 513586 708358
rect 513822 708122 549266 708358
rect 549502 708122 549586 708358
rect 549822 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect -5846 708090 589770 708122
rect -4886 707718 588810 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 23546 707718
rect 23782 707482 23866 707718
rect 24102 707482 59546 707718
rect 59782 707482 59866 707718
rect 60102 707482 95546 707718
rect 95782 707482 95866 707718
rect 96102 707482 131546 707718
rect 131782 707482 131866 707718
rect 132102 707482 167546 707718
rect 167782 707482 167866 707718
rect 168102 707482 203546 707718
rect 203782 707482 203866 707718
rect 204102 707482 239546 707718
rect 239782 707482 239866 707718
rect 240102 707482 275546 707718
rect 275782 707482 275866 707718
rect 276102 707482 311546 707718
rect 311782 707482 311866 707718
rect 312102 707482 347546 707718
rect 347782 707482 347866 707718
rect 348102 707482 383546 707718
rect 383782 707482 383866 707718
rect 384102 707482 419546 707718
rect 419782 707482 419866 707718
rect 420102 707482 455546 707718
rect 455782 707482 455866 707718
rect 456102 707482 491546 707718
rect 491782 707482 491866 707718
rect 492102 707482 527546 707718
rect 527782 707482 527866 707718
rect 528102 707482 563546 707718
rect 563782 707482 563866 707718
rect 564102 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect -4886 707398 588810 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 23546 707398
rect 23782 707162 23866 707398
rect 24102 707162 59546 707398
rect 59782 707162 59866 707398
rect 60102 707162 95546 707398
rect 95782 707162 95866 707398
rect 96102 707162 131546 707398
rect 131782 707162 131866 707398
rect 132102 707162 167546 707398
rect 167782 707162 167866 707398
rect 168102 707162 203546 707398
rect 203782 707162 203866 707398
rect 204102 707162 239546 707398
rect 239782 707162 239866 707398
rect 240102 707162 275546 707398
rect 275782 707162 275866 707398
rect 276102 707162 311546 707398
rect 311782 707162 311866 707398
rect 312102 707162 347546 707398
rect 347782 707162 347866 707398
rect 348102 707162 383546 707398
rect 383782 707162 383866 707398
rect 384102 707162 419546 707398
rect 419782 707162 419866 707398
rect 420102 707162 455546 707398
rect 455782 707162 455866 707398
rect 456102 707162 491546 707398
rect 491782 707162 491866 707398
rect 492102 707162 527546 707398
rect 527782 707162 527866 707398
rect 528102 707162 563546 707398
rect 563782 707162 563866 707398
rect 564102 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect -4886 707130 588810 707162
rect -3926 706758 587850 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 5546 706758
rect 5782 706522 5866 706758
rect 6102 706522 41546 706758
rect 41782 706522 41866 706758
rect 42102 706522 77546 706758
rect 77782 706522 77866 706758
rect 78102 706522 113546 706758
rect 113782 706522 113866 706758
rect 114102 706522 149546 706758
rect 149782 706522 149866 706758
rect 150102 706522 185546 706758
rect 185782 706522 185866 706758
rect 186102 706522 221546 706758
rect 221782 706522 221866 706758
rect 222102 706522 257546 706758
rect 257782 706522 257866 706758
rect 258102 706522 293546 706758
rect 293782 706522 293866 706758
rect 294102 706522 329546 706758
rect 329782 706522 329866 706758
rect 330102 706522 365546 706758
rect 365782 706522 365866 706758
rect 366102 706522 401546 706758
rect 401782 706522 401866 706758
rect 402102 706522 437546 706758
rect 437782 706522 437866 706758
rect 438102 706522 473546 706758
rect 473782 706522 473866 706758
rect 474102 706522 509546 706758
rect 509782 706522 509866 706758
rect 510102 706522 545546 706758
rect 545782 706522 545866 706758
rect 546102 706522 581546 706758
rect 581782 706522 581866 706758
rect 582102 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect -3926 706438 587850 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 5546 706438
rect 5782 706202 5866 706438
rect 6102 706202 41546 706438
rect 41782 706202 41866 706438
rect 42102 706202 77546 706438
rect 77782 706202 77866 706438
rect 78102 706202 113546 706438
rect 113782 706202 113866 706438
rect 114102 706202 149546 706438
rect 149782 706202 149866 706438
rect 150102 706202 185546 706438
rect 185782 706202 185866 706438
rect 186102 706202 221546 706438
rect 221782 706202 221866 706438
rect 222102 706202 257546 706438
rect 257782 706202 257866 706438
rect 258102 706202 293546 706438
rect 293782 706202 293866 706438
rect 294102 706202 329546 706438
rect 329782 706202 329866 706438
rect 330102 706202 365546 706438
rect 365782 706202 365866 706438
rect 366102 706202 401546 706438
rect 401782 706202 401866 706438
rect 402102 706202 437546 706438
rect 437782 706202 437866 706438
rect 438102 706202 473546 706438
rect 473782 706202 473866 706438
rect 474102 706202 509546 706438
rect 509782 706202 509866 706438
rect 510102 706202 545546 706438
rect 545782 706202 545866 706438
rect 546102 706202 581546 706438
rect 581782 706202 581866 706438
rect 582102 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect -3926 706170 587850 706202
rect -2966 705798 586890 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 19826 705798
rect 20062 705562 20146 705798
rect 20382 705562 55826 705798
rect 56062 705562 56146 705798
rect 56382 705562 91826 705798
rect 92062 705562 92146 705798
rect 92382 705562 127826 705798
rect 128062 705562 128146 705798
rect 128382 705562 163826 705798
rect 164062 705562 164146 705798
rect 164382 705562 199826 705798
rect 200062 705562 200146 705798
rect 200382 705562 235826 705798
rect 236062 705562 236146 705798
rect 236382 705562 271826 705798
rect 272062 705562 272146 705798
rect 272382 705562 307826 705798
rect 308062 705562 308146 705798
rect 308382 705562 343826 705798
rect 344062 705562 344146 705798
rect 344382 705562 379826 705798
rect 380062 705562 380146 705798
rect 380382 705562 415826 705798
rect 416062 705562 416146 705798
rect 416382 705562 451826 705798
rect 452062 705562 452146 705798
rect 452382 705562 487826 705798
rect 488062 705562 488146 705798
rect 488382 705562 523826 705798
rect 524062 705562 524146 705798
rect 524382 705562 559826 705798
rect 560062 705562 560146 705798
rect 560382 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect -2966 705478 586890 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 19826 705478
rect 20062 705242 20146 705478
rect 20382 705242 55826 705478
rect 56062 705242 56146 705478
rect 56382 705242 91826 705478
rect 92062 705242 92146 705478
rect 92382 705242 127826 705478
rect 128062 705242 128146 705478
rect 128382 705242 163826 705478
rect 164062 705242 164146 705478
rect 164382 705242 199826 705478
rect 200062 705242 200146 705478
rect 200382 705242 235826 705478
rect 236062 705242 236146 705478
rect 236382 705242 271826 705478
rect 272062 705242 272146 705478
rect 272382 705242 307826 705478
rect 308062 705242 308146 705478
rect 308382 705242 343826 705478
rect 344062 705242 344146 705478
rect 344382 705242 379826 705478
rect 380062 705242 380146 705478
rect 380382 705242 415826 705478
rect 416062 705242 416146 705478
rect 416382 705242 451826 705478
rect 452062 705242 452146 705478
rect 452382 705242 487826 705478
rect 488062 705242 488146 705478
rect 488382 705242 523826 705478
rect 524062 705242 524146 705478
rect 524382 705242 559826 705478
rect 560062 705242 560146 705478
rect 560382 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect -2966 705210 586890 705242
rect -2006 704838 585930 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect -2006 704518 585930 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect -2006 704250 585930 704282
rect -8726 698614 592650 698646
rect -8726 698378 -7734 698614
rect -7498 698378 -7414 698614
rect -7178 698378 12986 698614
rect 13222 698378 13306 698614
rect 13542 698378 48986 698614
rect 49222 698378 49306 698614
rect 49542 698378 84986 698614
rect 85222 698378 85306 698614
rect 85542 698378 120986 698614
rect 121222 698378 121306 698614
rect 121542 698378 156986 698614
rect 157222 698378 157306 698614
rect 157542 698378 192986 698614
rect 193222 698378 193306 698614
rect 193542 698378 228986 698614
rect 229222 698378 229306 698614
rect 229542 698378 264986 698614
rect 265222 698378 265306 698614
rect 265542 698378 300986 698614
rect 301222 698378 301306 698614
rect 301542 698378 336986 698614
rect 337222 698378 337306 698614
rect 337542 698378 372986 698614
rect 373222 698378 373306 698614
rect 373542 698378 408986 698614
rect 409222 698378 409306 698614
rect 409542 698378 444986 698614
rect 445222 698378 445306 698614
rect 445542 698378 480986 698614
rect 481222 698378 481306 698614
rect 481542 698378 516986 698614
rect 517222 698378 517306 698614
rect 517542 698378 552986 698614
rect 553222 698378 553306 698614
rect 553542 698378 591102 698614
rect 591338 698378 591422 698614
rect 591658 698378 592650 698614
rect -8726 698294 592650 698378
rect -8726 698058 -7734 698294
rect -7498 698058 -7414 698294
rect -7178 698058 12986 698294
rect 13222 698058 13306 698294
rect 13542 698058 48986 698294
rect 49222 698058 49306 698294
rect 49542 698058 84986 698294
rect 85222 698058 85306 698294
rect 85542 698058 120986 698294
rect 121222 698058 121306 698294
rect 121542 698058 156986 698294
rect 157222 698058 157306 698294
rect 157542 698058 192986 698294
rect 193222 698058 193306 698294
rect 193542 698058 228986 698294
rect 229222 698058 229306 698294
rect 229542 698058 264986 698294
rect 265222 698058 265306 698294
rect 265542 698058 300986 698294
rect 301222 698058 301306 698294
rect 301542 698058 336986 698294
rect 337222 698058 337306 698294
rect 337542 698058 372986 698294
rect 373222 698058 373306 698294
rect 373542 698058 408986 698294
rect 409222 698058 409306 698294
rect 409542 698058 444986 698294
rect 445222 698058 445306 698294
rect 445542 698058 480986 698294
rect 481222 698058 481306 698294
rect 481542 698058 516986 698294
rect 517222 698058 517306 698294
rect 517542 698058 552986 698294
rect 553222 698058 553306 698294
rect 553542 698058 591102 698294
rect 591338 698058 591422 698294
rect 591658 698058 592650 698294
rect -8726 698026 592650 698058
rect -6806 694894 590730 694926
rect -6806 694658 -5814 694894
rect -5578 694658 -5494 694894
rect -5258 694658 9266 694894
rect 9502 694658 9586 694894
rect 9822 694658 45266 694894
rect 45502 694658 45586 694894
rect 45822 694658 81266 694894
rect 81502 694658 81586 694894
rect 81822 694658 117266 694894
rect 117502 694658 117586 694894
rect 117822 694658 153266 694894
rect 153502 694658 153586 694894
rect 153822 694658 189266 694894
rect 189502 694658 189586 694894
rect 189822 694658 225266 694894
rect 225502 694658 225586 694894
rect 225822 694658 261266 694894
rect 261502 694658 261586 694894
rect 261822 694658 297266 694894
rect 297502 694658 297586 694894
rect 297822 694658 333266 694894
rect 333502 694658 333586 694894
rect 333822 694658 369266 694894
rect 369502 694658 369586 694894
rect 369822 694658 405266 694894
rect 405502 694658 405586 694894
rect 405822 694658 441266 694894
rect 441502 694658 441586 694894
rect 441822 694658 477266 694894
rect 477502 694658 477586 694894
rect 477822 694658 513266 694894
rect 513502 694658 513586 694894
rect 513822 694658 549266 694894
rect 549502 694658 549586 694894
rect 549822 694658 589182 694894
rect 589418 694658 589502 694894
rect 589738 694658 590730 694894
rect -6806 694574 590730 694658
rect -6806 694338 -5814 694574
rect -5578 694338 -5494 694574
rect -5258 694338 9266 694574
rect 9502 694338 9586 694574
rect 9822 694338 45266 694574
rect 45502 694338 45586 694574
rect 45822 694338 81266 694574
rect 81502 694338 81586 694574
rect 81822 694338 117266 694574
rect 117502 694338 117586 694574
rect 117822 694338 153266 694574
rect 153502 694338 153586 694574
rect 153822 694338 189266 694574
rect 189502 694338 189586 694574
rect 189822 694338 225266 694574
rect 225502 694338 225586 694574
rect 225822 694338 261266 694574
rect 261502 694338 261586 694574
rect 261822 694338 297266 694574
rect 297502 694338 297586 694574
rect 297822 694338 333266 694574
rect 333502 694338 333586 694574
rect 333822 694338 369266 694574
rect 369502 694338 369586 694574
rect 369822 694338 405266 694574
rect 405502 694338 405586 694574
rect 405822 694338 441266 694574
rect 441502 694338 441586 694574
rect 441822 694338 477266 694574
rect 477502 694338 477586 694574
rect 477822 694338 513266 694574
rect 513502 694338 513586 694574
rect 513822 694338 549266 694574
rect 549502 694338 549586 694574
rect 549822 694338 589182 694574
rect 589418 694338 589502 694574
rect 589738 694338 590730 694574
rect -6806 694306 590730 694338
rect -4886 691174 588810 691206
rect -4886 690938 -3894 691174
rect -3658 690938 -3574 691174
rect -3338 690938 5546 691174
rect 5782 690938 5866 691174
rect 6102 690938 41546 691174
rect 41782 690938 41866 691174
rect 42102 690938 77546 691174
rect 77782 690938 77866 691174
rect 78102 690938 113546 691174
rect 113782 690938 113866 691174
rect 114102 690938 149546 691174
rect 149782 690938 149866 691174
rect 150102 690938 185546 691174
rect 185782 690938 185866 691174
rect 186102 690938 221546 691174
rect 221782 690938 221866 691174
rect 222102 690938 257546 691174
rect 257782 690938 257866 691174
rect 258102 690938 293546 691174
rect 293782 690938 293866 691174
rect 294102 690938 329546 691174
rect 329782 690938 329866 691174
rect 330102 690938 365546 691174
rect 365782 690938 365866 691174
rect 366102 690938 401546 691174
rect 401782 690938 401866 691174
rect 402102 690938 437546 691174
rect 437782 690938 437866 691174
rect 438102 690938 473546 691174
rect 473782 690938 473866 691174
rect 474102 690938 509546 691174
rect 509782 690938 509866 691174
rect 510102 690938 545546 691174
rect 545782 690938 545866 691174
rect 546102 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 587262 691174
rect 587498 690938 587582 691174
rect 587818 690938 588810 691174
rect -4886 690854 588810 690938
rect -4886 690618 -3894 690854
rect -3658 690618 -3574 690854
rect -3338 690618 5546 690854
rect 5782 690618 5866 690854
rect 6102 690618 41546 690854
rect 41782 690618 41866 690854
rect 42102 690618 77546 690854
rect 77782 690618 77866 690854
rect 78102 690618 113546 690854
rect 113782 690618 113866 690854
rect 114102 690618 149546 690854
rect 149782 690618 149866 690854
rect 150102 690618 185546 690854
rect 185782 690618 185866 690854
rect 186102 690618 221546 690854
rect 221782 690618 221866 690854
rect 222102 690618 257546 690854
rect 257782 690618 257866 690854
rect 258102 690618 293546 690854
rect 293782 690618 293866 690854
rect 294102 690618 329546 690854
rect 329782 690618 329866 690854
rect 330102 690618 365546 690854
rect 365782 690618 365866 690854
rect 366102 690618 401546 690854
rect 401782 690618 401866 690854
rect 402102 690618 437546 690854
rect 437782 690618 437866 690854
rect 438102 690618 473546 690854
rect 473782 690618 473866 690854
rect 474102 690618 509546 690854
rect 509782 690618 509866 690854
rect 510102 690618 545546 690854
rect 545782 690618 545866 690854
rect 546102 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 587262 690854
rect 587498 690618 587582 690854
rect 587818 690618 588810 690854
rect -4886 690586 588810 690618
rect -2966 687454 586890 687486
rect -2966 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 586890 687454
rect -2966 687134 586890 687218
rect -2966 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 586890 687134
rect -2966 686866 586890 686898
rect -8726 680614 592650 680646
rect -8726 680378 -8694 680614
rect -8458 680378 -8374 680614
rect -8138 680378 30986 680614
rect 31222 680378 31306 680614
rect 31542 680378 66986 680614
rect 67222 680378 67306 680614
rect 67542 680378 102986 680614
rect 103222 680378 103306 680614
rect 103542 680378 138986 680614
rect 139222 680378 139306 680614
rect 139542 680378 174986 680614
rect 175222 680378 175306 680614
rect 175542 680378 210986 680614
rect 211222 680378 211306 680614
rect 211542 680378 246986 680614
rect 247222 680378 247306 680614
rect 247542 680378 282986 680614
rect 283222 680378 283306 680614
rect 283542 680378 318986 680614
rect 319222 680378 319306 680614
rect 319542 680378 354986 680614
rect 355222 680378 355306 680614
rect 355542 680378 390986 680614
rect 391222 680378 391306 680614
rect 391542 680378 426986 680614
rect 427222 680378 427306 680614
rect 427542 680378 462986 680614
rect 463222 680378 463306 680614
rect 463542 680378 498986 680614
rect 499222 680378 499306 680614
rect 499542 680378 534986 680614
rect 535222 680378 535306 680614
rect 535542 680378 570986 680614
rect 571222 680378 571306 680614
rect 571542 680378 592062 680614
rect 592298 680378 592382 680614
rect 592618 680378 592650 680614
rect -8726 680294 592650 680378
rect -8726 680058 -8694 680294
rect -8458 680058 -8374 680294
rect -8138 680058 30986 680294
rect 31222 680058 31306 680294
rect 31542 680058 66986 680294
rect 67222 680058 67306 680294
rect 67542 680058 102986 680294
rect 103222 680058 103306 680294
rect 103542 680058 138986 680294
rect 139222 680058 139306 680294
rect 139542 680058 174986 680294
rect 175222 680058 175306 680294
rect 175542 680058 210986 680294
rect 211222 680058 211306 680294
rect 211542 680058 246986 680294
rect 247222 680058 247306 680294
rect 247542 680058 282986 680294
rect 283222 680058 283306 680294
rect 283542 680058 318986 680294
rect 319222 680058 319306 680294
rect 319542 680058 354986 680294
rect 355222 680058 355306 680294
rect 355542 680058 390986 680294
rect 391222 680058 391306 680294
rect 391542 680058 426986 680294
rect 427222 680058 427306 680294
rect 427542 680058 462986 680294
rect 463222 680058 463306 680294
rect 463542 680058 498986 680294
rect 499222 680058 499306 680294
rect 499542 680058 534986 680294
rect 535222 680058 535306 680294
rect 535542 680058 570986 680294
rect 571222 680058 571306 680294
rect 571542 680058 592062 680294
rect 592298 680058 592382 680294
rect 592618 680058 592650 680294
rect -8726 680026 592650 680058
rect -6806 676894 590730 676926
rect -6806 676658 -6774 676894
rect -6538 676658 -6454 676894
rect -6218 676658 27266 676894
rect 27502 676658 27586 676894
rect 27822 676658 63266 676894
rect 63502 676658 63586 676894
rect 63822 676658 99266 676894
rect 99502 676658 99586 676894
rect 99822 676658 135266 676894
rect 135502 676658 135586 676894
rect 135822 676658 171266 676894
rect 171502 676658 171586 676894
rect 171822 676658 207266 676894
rect 207502 676658 207586 676894
rect 207822 676658 243266 676894
rect 243502 676658 243586 676894
rect 243822 676658 279266 676894
rect 279502 676658 279586 676894
rect 279822 676658 315266 676894
rect 315502 676658 315586 676894
rect 315822 676658 351266 676894
rect 351502 676658 351586 676894
rect 351822 676658 387266 676894
rect 387502 676658 387586 676894
rect 387822 676658 423266 676894
rect 423502 676658 423586 676894
rect 423822 676658 459266 676894
rect 459502 676658 459586 676894
rect 459822 676658 495266 676894
rect 495502 676658 495586 676894
rect 495822 676658 531266 676894
rect 531502 676658 531586 676894
rect 531822 676658 567266 676894
rect 567502 676658 567586 676894
rect 567822 676658 590142 676894
rect 590378 676658 590462 676894
rect 590698 676658 590730 676894
rect -6806 676574 590730 676658
rect -6806 676338 -6774 676574
rect -6538 676338 -6454 676574
rect -6218 676338 27266 676574
rect 27502 676338 27586 676574
rect 27822 676338 63266 676574
rect 63502 676338 63586 676574
rect 63822 676338 99266 676574
rect 99502 676338 99586 676574
rect 99822 676338 135266 676574
rect 135502 676338 135586 676574
rect 135822 676338 171266 676574
rect 171502 676338 171586 676574
rect 171822 676338 207266 676574
rect 207502 676338 207586 676574
rect 207822 676338 243266 676574
rect 243502 676338 243586 676574
rect 243822 676338 279266 676574
rect 279502 676338 279586 676574
rect 279822 676338 315266 676574
rect 315502 676338 315586 676574
rect 315822 676338 351266 676574
rect 351502 676338 351586 676574
rect 351822 676338 387266 676574
rect 387502 676338 387586 676574
rect 387822 676338 423266 676574
rect 423502 676338 423586 676574
rect 423822 676338 459266 676574
rect 459502 676338 459586 676574
rect 459822 676338 495266 676574
rect 495502 676338 495586 676574
rect 495822 676338 531266 676574
rect 531502 676338 531586 676574
rect 531822 676338 567266 676574
rect 567502 676338 567586 676574
rect 567822 676338 590142 676574
rect 590378 676338 590462 676574
rect 590698 676338 590730 676574
rect -6806 676306 590730 676338
rect -4886 673174 588810 673206
rect -4886 672938 -4854 673174
rect -4618 672938 -4534 673174
rect -4298 672938 23546 673174
rect 23782 672938 23866 673174
rect 24102 672938 59546 673174
rect 59782 672938 59866 673174
rect 60102 672938 95546 673174
rect 95782 672938 95866 673174
rect 96102 672938 131546 673174
rect 131782 672938 131866 673174
rect 132102 672938 167546 673174
rect 167782 672938 167866 673174
rect 168102 672938 203546 673174
rect 203782 672938 203866 673174
rect 204102 672938 239546 673174
rect 239782 672938 239866 673174
rect 240102 672938 275546 673174
rect 275782 672938 275866 673174
rect 276102 672938 311546 673174
rect 311782 672938 311866 673174
rect 312102 672938 347546 673174
rect 347782 672938 347866 673174
rect 348102 672938 383546 673174
rect 383782 672938 383866 673174
rect 384102 672938 419546 673174
rect 419782 672938 419866 673174
rect 420102 672938 455546 673174
rect 455782 672938 455866 673174
rect 456102 672938 491546 673174
rect 491782 672938 491866 673174
rect 492102 672938 527546 673174
rect 527782 672938 527866 673174
rect 528102 672938 563546 673174
rect 563782 672938 563866 673174
rect 564102 672938 588222 673174
rect 588458 672938 588542 673174
rect 588778 672938 588810 673174
rect -4886 672854 588810 672938
rect -4886 672618 -4854 672854
rect -4618 672618 -4534 672854
rect -4298 672618 23546 672854
rect 23782 672618 23866 672854
rect 24102 672618 59546 672854
rect 59782 672618 59866 672854
rect 60102 672618 95546 672854
rect 95782 672618 95866 672854
rect 96102 672618 131546 672854
rect 131782 672618 131866 672854
rect 132102 672618 167546 672854
rect 167782 672618 167866 672854
rect 168102 672618 203546 672854
rect 203782 672618 203866 672854
rect 204102 672618 239546 672854
rect 239782 672618 239866 672854
rect 240102 672618 275546 672854
rect 275782 672618 275866 672854
rect 276102 672618 311546 672854
rect 311782 672618 311866 672854
rect 312102 672618 347546 672854
rect 347782 672618 347866 672854
rect 348102 672618 383546 672854
rect 383782 672618 383866 672854
rect 384102 672618 419546 672854
rect 419782 672618 419866 672854
rect 420102 672618 455546 672854
rect 455782 672618 455866 672854
rect 456102 672618 491546 672854
rect 491782 672618 491866 672854
rect 492102 672618 527546 672854
rect 527782 672618 527866 672854
rect 528102 672618 563546 672854
rect 563782 672618 563866 672854
rect 564102 672618 588222 672854
rect 588458 672618 588542 672854
rect 588778 672618 588810 672854
rect -4886 672586 588810 672618
rect -2966 669454 586890 669486
rect -2966 669218 -2934 669454
rect -2698 669218 -2614 669454
rect -2378 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 586302 669454
rect 586538 669218 586622 669454
rect 586858 669218 586890 669454
rect -2966 669134 586890 669218
rect -2966 668898 -2934 669134
rect -2698 668898 -2614 669134
rect -2378 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 586302 669134
rect 586538 668898 586622 669134
rect 586858 668898 586890 669134
rect -2966 668866 586890 668898
rect -8726 662614 592650 662646
rect -8726 662378 -7734 662614
rect -7498 662378 -7414 662614
rect -7178 662378 12986 662614
rect 13222 662378 13306 662614
rect 13542 662378 48986 662614
rect 49222 662378 49306 662614
rect 49542 662378 84986 662614
rect 85222 662378 85306 662614
rect 85542 662378 120986 662614
rect 121222 662378 121306 662614
rect 121542 662378 156986 662614
rect 157222 662378 157306 662614
rect 157542 662378 192986 662614
rect 193222 662378 193306 662614
rect 193542 662378 228986 662614
rect 229222 662378 229306 662614
rect 229542 662378 264986 662614
rect 265222 662378 265306 662614
rect 265542 662378 300986 662614
rect 301222 662378 301306 662614
rect 301542 662378 336986 662614
rect 337222 662378 337306 662614
rect 337542 662378 372986 662614
rect 373222 662378 373306 662614
rect 373542 662378 408986 662614
rect 409222 662378 409306 662614
rect 409542 662378 444986 662614
rect 445222 662378 445306 662614
rect 445542 662378 480986 662614
rect 481222 662378 481306 662614
rect 481542 662378 516986 662614
rect 517222 662378 517306 662614
rect 517542 662378 552986 662614
rect 553222 662378 553306 662614
rect 553542 662378 591102 662614
rect 591338 662378 591422 662614
rect 591658 662378 592650 662614
rect -8726 662294 592650 662378
rect -8726 662058 -7734 662294
rect -7498 662058 -7414 662294
rect -7178 662058 12986 662294
rect 13222 662058 13306 662294
rect 13542 662058 48986 662294
rect 49222 662058 49306 662294
rect 49542 662058 84986 662294
rect 85222 662058 85306 662294
rect 85542 662058 120986 662294
rect 121222 662058 121306 662294
rect 121542 662058 156986 662294
rect 157222 662058 157306 662294
rect 157542 662058 192986 662294
rect 193222 662058 193306 662294
rect 193542 662058 228986 662294
rect 229222 662058 229306 662294
rect 229542 662058 264986 662294
rect 265222 662058 265306 662294
rect 265542 662058 300986 662294
rect 301222 662058 301306 662294
rect 301542 662058 336986 662294
rect 337222 662058 337306 662294
rect 337542 662058 372986 662294
rect 373222 662058 373306 662294
rect 373542 662058 408986 662294
rect 409222 662058 409306 662294
rect 409542 662058 444986 662294
rect 445222 662058 445306 662294
rect 445542 662058 480986 662294
rect 481222 662058 481306 662294
rect 481542 662058 516986 662294
rect 517222 662058 517306 662294
rect 517542 662058 552986 662294
rect 553222 662058 553306 662294
rect 553542 662058 591102 662294
rect 591338 662058 591422 662294
rect 591658 662058 592650 662294
rect -8726 662026 592650 662058
rect -6806 658894 590730 658926
rect -6806 658658 -5814 658894
rect -5578 658658 -5494 658894
rect -5258 658658 9266 658894
rect 9502 658658 9586 658894
rect 9822 658658 45266 658894
rect 45502 658658 45586 658894
rect 45822 658658 81266 658894
rect 81502 658658 81586 658894
rect 81822 658658 117266 658894
rect 117502 658658 117586 658894
rect 117822 658658 153266 658894
rect 153502 658658 153586 658894
rect 153822 658658 189266 658894
rect 189502 658658 189586 658894
rect 189822 658658 225266 658894
rect 225502 658658 225586 658894
rect 225822 658658 261266 658894
rect 261502 658658 261586 658894
rect 261822 658658 297266 658894
rect 297502 658658 297586 658894
rect 297822 658658 333266 658894
rect 333502 658658 333586 658894
rect 333822 658658 369266 658894
rect 369502 658658 369586 658894
rect 369822 658658 405266 658894
rect 405502 658658 405586 658894
rect 405822 658658 441266 658894
rect 441502 658658 441586 658894
rect 441822 658658 477266 658894
rect 477502 658658 477586 658894
rect 477822 658658 513266 658894
rect 513502 658658 513586 658894
rect 513822 658658 549266 658894
rect 549502 658658 549586 658894
rect 549822 658658 589182 658894
rect 589418 658658 589502 658894
rect 589738 658658 590730 658894
rect -6806 658574 590730 658658
rect -6806 658338 -5814 658574
rect -5578 658338 -5494 658574
rect -5258 658338 9266 658574
rect 9502 658338 9586 658574
rect 9822 658338 45266 658574
rect 45502 658338 45586 658574
rect 45822 658338 81266 658574
rect 81502 658338 81586 658574
rect 81822 658338 117266 658574
rect 117502 658338 117586 658574
rect 117822 658338 153266 658574
rect 153502 658338 153586 658574
rect 153822 658338 189266 658574
rect 189502 658338 189586 658574
rect 189822 658338 225266 658574
rect 225502 658338 225586 658574
rect 225822 658338 261266 658574
rect 261502 658338 261586 658574
rect 261822 658338 297266 658574
rect 297502 658338 297586 658574
rect 297822 658338 333266 658574
rect 333502 658338 333586 658574
rect 333822 658338 369266 658574
rect 369502 658338 369586 658574
rect 369822 658338 405266 658574
rect 405502 658338 405586 658574
rect 405822 658338 441266 658574
rect 441502 658338 441586 658574
rect 441822 658338 477266 658574
rect 477502 658338 477586 658574
rect 477822 658338 513266 658574
rect 513502 658338 513586 658574
rect 513822 658338 549266 658574
rect 549502 658338 549586 658574
rect 549822 658338 589182 658574
rect 589418 658338 589502 658574
rect 589738 658338 590730 658574
rect -6806 658306 590730 658338
rect -4886 655174 588810 655206
rect -4886 654938 -3894 655174
rect -3658 654938 -3574 655174
rect -3338 654938 5546 655174
rect 5782 654938 5866 655174
rect 6102 654938 41546 655174
rect 41782 654938 41866 655174
rect 42102 654938 77546 655174
rect 77782 654938 77866 655174
rect 78102 654938 113546 655174
rect 113782 654938 113866 655174
rect 114102 654938 149546 655174
rect 149782 654938 149866 655174
rect 150102 654938 185546 655174
rect 185782 654938 185866 655174
rect 186102 654938 221546 655174
rect 221782 654938 221866 655174
rect 222102 654938 257546 655174
rect 257782 654938 257866 655174
rect 258102 654938 293546 655174
rect 293782 654938 293866 655174
rect 294102 654938 329546 655174
rect 329782 654938 329866 655174
rect 330102 654938 365546 655174
rect 365782 654938 365866 655174
rect 366102 654938 401546 655174
rect 401782 654938 401866 655174
rect 402102 654938 437546 655174
rect 437782 654938 437866 655174
rect 438102 654938 473546 655174
rect 473782 654938 473866 655174
rect 474102 654938 509546 655174
rect 509782 654938 509866 655174
rect 510102 654938 545546 655174
rect 545782 654938 545866 655174
rect 546102 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 587262 655174
rect 587498 654938 587582 655174
rect 587818 654938 588810 655174
rect -4886 654854 588810 654938
rect -4886 654618 -3894 654854
rect -3658 654618 -3574 654854
rect -3338 654618 5546 654854
rect 5782 654618 5866 654854
rect 6102 654618 41546 654854
rect 41782 654618 41866 654854
rect 42102 654618 77546 654854
rect 77782 654618 77866 654854
rect 78102 654618 113546 654854
rect 113782 654618 113866 654854
rect 114102 654618 149546 654854
rect 149782 654618 149866 654854
rect 150102 654618 185546 654854
rect 185782 654618 185866 654854
rect 186102 654618 221546 654854
rect 221782 654618 221866 654854
rect 222102 654618 257546 654854
rect 257782 654618 257866 654854
rect 258102 654618 293546 654854
rect 293782 654618 293866 654854
rect 294102 654618 329546 654854
rect 329782 654618 329866 654854
rect 330102 654618 365546 654854
rect 365782 654618 365866 654854
rect 366102 654618 401546 654854
rect 401782 654618 401866 654854
rect 402102 654618 437546 654854
rect 437782 654618 437866 654854
rect 438102 654618 473546 654854
rect 473782 654618 473866 654854
rect 474102 654618 509546 654854
rect 509782 654618 509866 654854
rect 510102 654618 545546 654854
rect 545782 654618 545866 654854
rect 546102 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 587262 654854
rect 587498 654618 587582 654854
rect 587818 654618 588810 654854
rect -4886 654586 588810 654618
rect -2966 651454 586890 651486
rect -2966 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 586890 651454
rect -2966 651134 586890 651218
rect -2966 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 586890 651134
rect -2966 650866 586890 650898
rect -8726 644614 592650 644646
rect -8726 644378 -8694 644614
rect -8458 644378 -8374 644614
rect -8138 644378 30986 644614
rect 31222 644378 31306 644614
rect 31542 644378 66986 644614
rect 67222 644378 67306 644614
rect 67542 644378 102986 644614
rect 103222 644378 103306 644614
rect 103542 644378 138986 644614
rect 139222 644378 139306 644614
rect 139542 644378 174986 644614
rect 175222 644378 175306 644614
rect 175542 644378 210986 644614
rect 211222 644378 211306 644614
rect 211542 644378 246986 644614
rect 247222 644378 247306 644614
rect 247542 644378 282986 644614
rect 283222 644378 283306 644614
rect 283542 644378 318986 644614
rect 319222 644378 319306 644614
rect 319542 644378 354986 644614
rect 355222 644378 355306 644614
rect 355542 644378 390986 644614
rect 391222 644378 391306 644614
rect 391542 644378 426986 644614
rect 427222 644378 427306 644614
rect 427542 644378 462986 644614
rect 463222 644378 463306 644614
rect 463542 644378 498986 644614
rect 499222 644378 499306 644614
rect 499542 644378 534986 644614
rect 535222 644378 535306 644614
rect 535542 644378 570986 644614
rect 571222 644378 571306 644614
rect 571542 644378 592062 644614
rect 592298 644378 592382 644614
rect 592618 644378 592650 644614
rect -8726 644294 592650 644378
rect -8726 644058 -8694 644294
rect -8458 644058 -8374 644294
rect -8138 644058 30986 644294
rect 31222 644058 31306 644294
rect 31542 644058 66986 644294
rect 67222 644058 67306 644294
rect 67542 644058 102986 644294
rect 103222 644058 103306 644294
rect 103542 644058 138986 644294
rect 139222 644058 139306 644294
rect 139542 644058 174986 644294
rect 175222 644058 175306 644294
rect 175542 644058 210986 644294
rect 211222 644058 211306 644294
rect 211542 644058 246986 644294
rect 247222 644058 247306 644294
rect 247542 644058 282986 644294
rect 283222 644058 283306 644294
rect 283542 644058 318986 644294
rect 319222 644058 319306 644294
rect 319542 644058 354986 644294
rect 355222 644058 355306 644294
rect 355542 644058 390986 644294
rect 391222 644058 391306 644294
rect 391542 644058 426986 644294
rect 427222 644058 427306 644294
rect 427542 644058 462986 644294
rect 463222 644058 463306 644294
rect 463542 644058 498986 644294
rect 499222 644058 499306 644294
rect 499542 644058 534986 644294
rect 535222 644058 535306 644294
rect 535542 644058 570986 644294
rect 571222 644058 571306 644294
rect 571542 644058 592062 644294
rect 592298 644058 592382 644294
rect 592618 644058 592650 644294
rect -8726 644026 592650 644058
rect -6806 640894 590730 640926
rect -6806 640658 -6774 640894
rect -6538 640658 -6454 640894
rect -6218 640658 27266 640894
rect 27502 640658 27586 640894
rect 27822 640658 63266 640894
rect 63502 640658 63586 640894
rect 63822 640658 99266 640894
rect 99502 640658 99586 640894
rect 99822 640658 135266 640894
rect 135502 640658 135586 640894
rect 135822 640658 171266 640894
rect 171502 640658 171586 640894
rect 171822 640658 207266 640894
rect 207502 640658 207586 640894
rect 207822 640658 243266 640894
rect 243502 640658 243586 640894
rect 243822 640658 279266 640894
rect 279502 640658 279586 640894
rect 279822 640658 315266 640894
rect 315502 640658 315586 640894
rect 315822 640658 351266 640894
rect 351502 640658 351586 640894
rect 351822 640658 387266 640894
rect 387502 640658 387586 640894
rect 387822 640658 423266 640894
rect 423502 640658 423586 640894
rect 423822 640658 459266 640894
rect 459502 640658 459586 640894
rect 459822 640658 495266 640894
rect 495502 640658 495586 640894
rect 495822 640658 531266 640894
rect 531502 640658 531586 640894
rect 531822 640658 567266 640894
rect 567502 640658 567586 640894
rect 567822 640658 590142 640894
rect 590378 640658 590462 640894
rect 590698 640658 590730 640894
rect -6806 640574 590730 640658
rect -6806 640338 -6774 640574
rect -6538 640338 -6454 640574
rect -6218 640338 27266 640574
rect 27502 640338 27586 640574
rect 27822 640338 63266 640574
rect 63502 640338 63586 640574
rect 63822 640338 99266 640574
rect 99502 640338 99586 640574
rect 99822 640338 135266 640574
rect 135502 640338 135586 640574
rect 135822 640338 171266 640574
rect 171502 640338 171586 640574
rect 171822 640338 207266 640574
rect 207502 640338 207586 640574
rect 207822 640338 243266 640574
rect 243502 640338 243586 640574
rect 243822 640338 279266 640574
rect 279502 640338 279586 640574
rect 279822 640338 315266 640574
rect 315502 640338 315586 640574
rect 315822 640338 351266 640574
rect 351502 640338 351586 640574
rect 351822 640338 387266 640574
rect 387502 640338 387586 640574
rect 387822 640338 423266 640574
rect 423502 640338 423586 640574
rect 423822 640338 459266 640574
rect 459502 640338 459586 640574
rect 459822 640338 495266 640574
rect 495502 640338 495586 640574
rect 495822 640338 531266 640574
rect 531502 640338 531586 640574
rect 531822 640338 567266 640574
rect 567502 640338 567586 640574
rect 567822 640338 590142 640574
rect 590378 640338 590462 640574
rect 590698 640338 590730 640574
rect -6806 640306 590730 640338
rect -4886 637174 588810 637206
rect -4886 636938 -4854 637174
rect -4618 636938 -4534 637174
rect -4298 636938 23546 637174
rect 23782 636938 23866 637174
rect 24102 636938 59546 637174
rect 59782 636938 59866 637174
rect 60102 636938 95546 637174
rect 95782 636938 95866 637174
rect 96102 636938 131546 637174
rect 131782 636938 131866 637174
rect 132102 636938 167546 637174
rect 167782 636938 167866 637174
rect 168102 636938 203546 637174
rect 203782 636938 203866 637174
rect 204102 636938 239546 637174
rect 239782 636938 239866 637174
rect 240102 636938 275546 637174
rect 275782 636938 275866 637174
rect 276102 636938 311546 637174
rect 311782 636938 311866 637174
rect 312102 636938 347546 637174
rect 347782 636938 347866 637174
rect 348102 636938 383546 637174
rect 383782 636938 383866 637174
rect 384102 636938 419546 637174
rect 419782 636938 419866 637174
rect 420102 636938 455546 637174
rect 455782 636938 455866 637174
rect 456102 636938 491546 637174
rect 491782 636938 491866 637174
rect 492102 636938 527546 637174
rect 527782 636938 527866 637174
rect 528102 636938 563546 637174
rect 563782 636938 563866 637174
rect 564102 636938 588222 637174
rect 588458 636938 588542 637174
rect 588778 636938 588810 637174
rect -4886 636854 588810 636938
rect -4886 636618 -4854 636854
rect -4618 636618 -4534 636854
rect -4298 636618 23546 636854
rect 23782 636618 23866 636854
rect 24102 636618 59546 636854
rect 59782 636618 59866 636854
rect 60102 636618 95546 636854
rect 95782 636618 95866 636854
rect 96102 636618 131546 636854
rect 131782 636618 131866 636854
rect 132102 636618 167546 636854
rect 167782 636618 167866 636854
rect 168102 636618 203546 636854
rect 203782 636618 203866 636854
rect 204102 636618 239546 636854
rect 239782 636618 239866 636854
rect 240102 636618 275546 636854
rect 275782 636618 275866 636854
rect 276102 636618 311546 636854
rect 311782 636618 311866 636854
rect 312102 636618 347546 636854
rect 347782 636618 347866 636854
rect 348102 636618 383546 636854
rect 383782 636618 383866 636854
rect 384102 636618 419546 636854
rect 419782 636618 419866 636854
rect 420102 636618 455546 636854
rect 455782 636618 455866 636854
rect 456102 636618 491546 636854
rect 491782 636618 491866 636854
rect 492102 636618 527546 636854
rect 527782 636618 527866 636854
rect 528102 636618 563546 636854
rect 563782 636618 563866 636854
rect 564102 636618 588222 636854
rect 588458 636618 588542 636854
rect 588778 636618 588810 636854
rect -4886 636586 588810 636618
rect -2966 633454 586890 633486
rect -2966 633218 -2934 633454
rect -2698 633218 -2614 633454
rect -2378 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 586302 633454
rect 586538 633218 586622 633454
rect 586858 633218 586890 633454
rect -2966 633134 586890 633218
rect -2966 632898 -2934 633134
rect -2698 632898 -2614 633134
rect -2378 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 586302 633134
rect 586538 632898 586622 633134
rect 586858 632898 586890 633134
rect -2966 632866 586890 632898
rect -8726 626614 592650 626646
rect -8726 626378 -7734 626614
rect -7498 626378 -7414 626614
rect -7178 626378 12986 626614
rect 13222 626378 13306 626614
rect 13542 626378 48986 626614
rect 49222 626378 49306 626614
rect 49542 626378 84986 626614
rect 85222 626378 85306 626614
rect 85542 626378 120986 626614
rect 121222 626378 121306 626614
rect 121542 626378 156986 626614
rect 157222 626378 157306 626614
rect 157542 626378 192986 626614
rect 193222 626378 193306 626614
rect 193542 626378 228986 626614
rect 229222 626378 229306 626614
rect 229542 626378 264986 626614
rect 265222 626378 265306 626614
rect 265542 626378 300986 626614
rect 301222 626378 301306 626614
rect 301542 626378 336986 626614
rect 337222 626378 337306 626614
rect 337542 626378 372986 626614
rect 373222 626378 373306 626614
rect 373542 626378 408986 626614
rect 409222 626378 409306 626614
rect 409542 626378 444986 626614
rect 445222 626378 445306 626614
rect 445542 626378 480986 626614
rect 481222 626378 481306 626614
rect 481542 626378 516986 626614
rect 517222 626378 517306 626614
rect 517542 626378 552986 626614
rect 553222 626378 553306 626614
rect 553542 626378 591102 626614
rect 591338 626378 591422 626614
rect 591658 626378 592650 626614
rect -8726 626294 592650 626378
rect -8726 626058 -7734 626294
rect -7498 626058 -7414 626294
rect -7178 626058 12986 626294
rect 13222 626058 13306 626294
rect 13542 626058 48986 626294
rect 49222 626058 49306 626294
rect 49542 626058 84986 626294
rect 85222 626058 85306 626294
rect 85542 626058 120986 626294
rect 121222 626058 121306 626294
rect 121542 626058 156986 626294
rect 157222 626058 157306 626294
rect 157542 626058 192986 626294
rect 193222 626058 193306 626294
rect 193542 626058 228986 626294
rect 229222 626058 229306 626294
rect 229542 626058 264986 626294
rect 265222 626058 265306 626294
rect 265542 626058 300986 626294
rect 301222 626058 301306 626294
rect 301542 626058 336986 626294
rect 337222 626058 337306 626294
rect 337542 626058 372986 626294
rect 373222 626058 373306 626294
rect 373542 626058 408986 626294
rect 409222 626058 409306 626294
rect 409542 626058 444986 626294
rect 445222 626058 445306 626294
rect 445542 626058 480986 626294
rect 481222 626058 481306 626294
rect 481542 626058 516986 626294
rect 517222 626058 517306 626294
rect 517542 626058 552986 626294
rect 553222 626058 553306 626294
rect 553542 626058 591102 626294
rect 591338 626058 591422 626294
rect 591658 626058 592650 626294
rect -8726 626026 592650 626058
rect -6806 622894 590730 622926
rect -6806 622658 -5814 622894
rect -5578 622658 -5494 622894
rect -5258 622658 9266 622894
rect 9502 622658 9586 622894
rect 9822 622658 45266 622894
rect 45502 622658 45586 622894
rect 45822 622658 81266 622894
rect 81502 622658 81586 622894
rect 81822 622658 117266 622894
rect 117502 622658 117586 622894
rect 117822 622658 153266 622894
rect 153502 622658 153586 622894
rect 153822 622658 189266 622894
rect 189502 622658 189586 622894
rect 189822 622658 225266 622894
rect 225502 622658 225586 622894
rect 225822 622658 261266 622894
rect 261502 622658 261586 622894
rect 261822 622658 297266 622894
rect 297502 622658 297586 622894
rect 297822 622658 333266 622894
rect 333502 622658 333586 622894
rect 333822 622658 369266 622894
rect 369502 622658 369586 622894
rect 369822 622658 405266 622894
rect 405502 622658 405586 622894
rect 405822 622658 441266 622894
rect 441502 622658 441586 622894
rect 441822 622658 477266 622894
rect 477502 622658 477586 622894
rect 477822 622658 513266 622894
rect 513502 622658 513586 622894
rect 513822 622658 549266 622894
rect 549502 622658 549586 622894
rect 549822 622658 589182 622894
rect 589418 622658 589502 622894
rect 589738 622658 590730 622894
rect -6806 622574 590730 622658
rect -6806 622338 -5814 622574
rect -5578 622338 -5494 622574
rect -5258 622338 9266 622574
rect 9502 622338 9586 622574
rect 9822 622338 45266 622574
rect 45502 622338 45586 622574
rect 45822 622338 81266 622574
rect 81502 622338 81586 622574
rect 81822 622338 117266 622574
rect 117502 622338 117586 622574
rect 117822 622338 153266 622574
rect 153502 622338 153586 622574
rect 153822 622338 189266 622574
rect 189502 622338 189586 622574
rect 189822 622338 225266 622574
rect 225502 622338 225586 622574
rect 225822 622338 261266 622574
rect 261502 622338 261586 622574
rect 261822 622338 297266 622574
rect 297502 622338 297586 622574
rect 297822 622338 333266 622574
rect 333502 622338 333586 622574
rect 333822 622338 369266 622574
rect 369502 622338 369586 622574
rect 369822 622338 405266 622574
rect 405502 622338 405586 622574
rect 405822 622338 441266 622574
rect 441502 622338 441586 622574
rect 441822 622338 477266 622574
rect 477502 622338 477586 622574
rect 477822 622338 513266 622574
rect 513502 622338 513586 622574
rect 513822 622338 549266 622574
rect 549502 622338 549586 622574
rect 549822 622338 589182 622574
rect 589418 622338 589502 622574
rect 589738 622338 590730 622574
rect -6806 622306 590730 622338
rect -4886 619174 588810 619206
rect -4886 618938 -3894 619174
rect -3658 618938 -3574 619174
rect -3338 618938 5546 619174
rect 5782 618938 5866 619174
rect 6102 618938 41546 619174
rect 41782 618938 41866 619174
rect 42102 618938 77546 619174
rect 77782 618938 77866 619174
rect 78102 618938 113546 619174
rect 113782 618938 113866 619174
rect 114102 618938 149546 619174
rect 149782 618938 149866 619174
rect 150102 618938 185546 619174
rect 185782 618938 185866 619174
rect 186102 618938 221546 619174
rect 221782 618938 221866 619174
rect 222102 618938 257546 619174
rect 257782 618938 257866 619174
rect 258102 618938 293546 619174
rect 293782 618938 293866 619174
rect 294102 618938 329546 619174
rect 329782 618938 329866 619174
rect 330102 618938 365546 619174
rect 365782 618938 365866 619174
rect 366102 618938 401546 619174
rect 401782 618938 401866 619174
rect 402102 618938 437546 619174
rect 437782 618938 437866 619174
rect 438102 618938 473546 619174
rect 473782 618938 473866 619174
rect 474102 618938 509546 619174
rect 509782 618938 509866 619174
rect 510102 618938 545546 619174
rect 545782 618938 545866 619174
rect 546102 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 587262 619174
rect 587498 618938 587582 619174
rect 587818 618938 588810 619174
rect -4886 618854 588810 618938
rect -4886 618618 -3894 618854
rect -3658 618618 -3574 618854
rect -3338 618618 5546 618854
rect 5782 618618 5866 618854
rect 6102 618618 41546 618854
rect 41782 618618 41866 618854
rect 42102 618618 77546 618854
rect 77782 618618 77866 618854
rect 78102 618618 113546 618854
rect 113782 618618 113866 618854
rect 114102 618618 149546 618854
rect 149782 618618 149866 618854
rect 150102 618618 185546 618854
rect 185782 618618 185866 618854
rect 186102 618618 221546 618854
rect 221782 618618 221866 618854
rect 222102 618618 257546 618854
rect 257782 618618 257866 618854
rect 258102 618618 293546 618854
rect 293782 618618 293866 618854
rect 294102 618618 329546 618854
rect 329782 618618 329866 618854
rect 330102 618618 365546 618854
rect 365782 618618 365866 618854
rect 366102 618618 401546 618854
rect 401782 618618 401866 618854
rect 402102 618618 437546 618854
rect 437782 618618 437866 618854
rect 438102 618618 473546 618854
rect 473782 618618 473866 618854
rect 474102 618618 509546 618854
rect 509782 618618 509866 618854
rect 510102 618618 545546 618854
rect 545782 618618 545866 618854
rect 546102 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 587262 618854
rect 587498 618618 587582 618854
rect 587818 618618 588810 618854
rect -4886 618586 588810 618618
rect -2966 615454 586890 615486
rect -2966 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 586890 615454
rect -2966 615134 586890 615218
rect -2966 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 586890 615134
rect -2966 614866 586890 614898
rect -8726 608614 592650 608646
rect -8726 608378 -8694 608614
rect -8458 608378 -8374 608614
rect -8138 608378 30986 608614
rect 31222 608378 31306 608614
rect 31542 608378 66986 608614
rect 67222 608378 67306 608614
rect 67542 608378 102986 608614
rect 103222 608378 103306 608614
rect 103542 608378 138986 608614
rect 139222 608378 139306 608614
rect 139542 608378 174986 608614
rect 175222 608378 175306 608614
rect 175542 608378 210986 608614
rect 211222 608378 211306 608614
rect 211542 608378 246986 608614
rect 247222 608378 247306 608614
rect 247542 608378 282986 608614
rect 283222 608378 283306 608614
rect 283542 608378 318986 608614
rect 319222 608378 319306 608614
rect 319542 608378 354986 608614
rect 355222 608378 355306 608614
rect 355542 608378 390986 608614
rect 391222 608378 391306 608614
rect 391542 608378 426986 608614
rect 427222 608378 427306 608614
rect 427542 608378 462986 608614
rect 463222 608378 463306 608614
rect 463542 608378 498986 608614
rect 499222 608378 499306 608614
rect 499542 608378 534986 608614
rect 535222 608378 535306 608614
rect 535542 608378 570986 608614
rect 571222 608378 571306 608614
rect 571542 608378 592062 608614
rect 592298 608378 592382 608614
rect 592618 608378 592650 608614
rect -8726 608294 592650 608378
rect -8726 608058 -8694 608294
rect -8458 608058 -8374 608294
rect -8138 608058 30986 608294
rect 31222 608058 31306 608294
rect 31542 608058 66986 608294
rect 67222 608058 67306 608294
rect 67542 608058 102986 608294
rect 103222 608058 103306 608294
rect 103542 608058 138986 608294
rect 139222 608058 139306 608294
rect 139542 608058 174986 608294
rect 175222 608058 175306 608294
rect 175542 608058 210986 608294
rect 211222 608058 211306 608294
rect 211542 608058 246986 608294
rect 247222 608058 247306 608294
rect 247542 608058 282986 608294
rect 283222 608058 283306 608294
rect 283542 608058 318986 608294
rect 319222 608058 319306 608294
rect 319542 608058 354986 608294
rect 355222 608058 355306 608294
rect 355542 608058 390986 608294
rect 391222 608058 391306 608294
rect 391542 608058 426986 608294
rect 427222 608058 427306 608294
rect 427542 608058 462986 608294
rect 463222 608058 463306 608294
rect 463542 608058 498986 608294
rect 499222 608058 499306 608294
rect 499542 608058 534986 608294
rect 535222 608058 535306 608294
rect 535542 608058 570986 608294
rect 571222 608058 571306 608294
rect 571542 608058 592062 608294
rect 592298 608058 592382 608294
rect 592618 608058 592650 608294
rect -8726 608026 592650 608058
rect -6806 604894 590730 604926
rect -6806 604658 -6774 604894
rect -6538 604658 -6454 604894
rect -6218 604658 27266 604894
rect 27502 604658 27586 604894
rect 27822 604658 63266 604894
rect 63502 604658 63586 604894
rect 63822 604658 99266 604894
rect 99502 604658 99586 604894
rect 99822 604658 135266 604894
rect 135502 604658 135586 604894
rect 135822 604658 171266 604894
rect 171502 604658 171586 604894
rect 171822 604658 207266 604894
rect 207502 604658 207586 604894
rect 207822 604658 243266 604894
rect 243502 604658 243586 604894
rect 243822 604658 279266 604894
rect 279502 604658 279586 604894
rect 279822 604658 315266 604894
rect 315502 604658 315586 604894
rect 315822 604658 351266 604894
rect 351502 604658 351586 604894
rect 351822 604658 387266 604894
rect 387502 604658 387586 604894
rect 387822 604658 423266 604894
rect 423502 604658 423586 604894
rect 423822 604658 459266 604894
rect 459502 604658 459586 604894
rect 459822 604658 495266 604894
rect 495502 604658 495586 604894
rect 495822 604658 531266 604894
rect 531502 604658 531586 604894
rect 531822 604658 567266 604894
rect 567502 604658 567586 604894
rect 567822 604658 590142 604894
rect 590378 604658 590462 604894
rect 590698 604658 590730 604894
rect -6806 604574 590730 604658
rect -6806 604338 -6774 604574
rect -6538 604338 -6454 604574
rect -6218 604338 27266 604574
rect 27502 604338 27586 604574
rect 27822 604338 63266 604574
rect 63502 604338 63586 604574
rect 63822 604338 99266 604574
rect 99502 604338 99586 604574
rect 99822 604338 135266 604574
rect 135502 604338 135586 604574
rect 135822 604338 171266 604574
rect 171502 604338 171586 604574
rect 171822 604338 207266 604574
rect 207502 604338 207586 604574
rect 207822 604338 243266 604574
rect 243502 604338 243586 604574
rect 243822 604338 279266 604574
rect 279502 604338 279586 604574
rect 279822 604338 315266 604574
rect 315502 604338 315586 604574
rect 315822 604338 351266 604574
rect 351502 604338 351586 604574
rect 351822 604338 387266 604574
rect 387502 604338 387586 604574
rect 387822 604338 423266 604574
rect 423502 604338 423586 604574
rect 423822 604338 459266 604574
rect 459502 604338 459586 604574
rect 459822 604338 495266 604574
rect 495502 604338 495586 604574
rect 495822 604338 531266 604574
rect 531502 604338 531586 604574
rect 531822 604338 567266 604574
rect 567502 604338 567586 604574
rect 567822 604338 590142 604574
rect 590378 604338 590462 604574
rect 590698 604338 590730 604574
rect -6806 604306 590730 604338
rect -4886 601174 588810 601206
rect -4886 600938 -4854 601174
rect -4618 600938 -4534 601174
rect -4298 600938 23546 601174
rect 23782 600938 23866 601174
rect 24102 600938 59546 601174
rect 59782 600938 59866 601174
rect 60102 600938 95546 601174
rect 95782 600938 95866 601174
rect 96102 600938 131546 601174
rect 131782 600938 131866 601174
rect 132102 600938 167546 601174
rect 167782 600938 167866 601174
rect 168102 600938 203546 601174
rect 203782 600938 203866 601174
rect 204102 600938 239546 601174
rect 239782 600938 239866 601174
rect 240102 600938 275546 601174
rect 275782 600938 275866 601174
rect 276102 600938 311546 601174
rect 311782 600938 311866 601174
rect 312102 600938 347546 601174
rect 347782 600938 347866 601174
rect 348102 600938 383546 601174
rect 383782 600938 383866 601174
rect 384102 600938 419546 601174
rect 419782 600938 419866 601174
rect 420102 600938 455546 601174
rect 455782 600938 455866 601174
rect 456102 600938 491546 601174
rect 491782 600938 491866 601174
rect 492102 600938 527546 601174
rect 527782 600938 527866 601174
rect 528102 600938 563546 601174
rect 563782 600938 563866 601174
rect 564102 600938 588222 601174
rect 588458 600938 588542 601174
rect 588778 600938 588810 601174
rect -4886 600854 588810 600938
rect -4886 600618 -4854 600854
rect -4618 600618 -4534 600854
rect -4298 600618 23546 600854
rect 23782 600618 23866 600854
rect 24102 600618 59546 600854
rect 59782 600618 59866 600854
rect 60102 600618 95546 600854
rect 95782 600618 95866 600854
rect 96102 600618 131546 600854
rect 131782 600618 131866 600854
rect 132102 600618 167546 600854
rect 167782 600618 167866 600854
rect 168102 600618 203546 600854
rect 203782 600618 203866 600854
rect 204102 600618 239546 600854
rect 239782 600618 239866 600854
rect 240102 600618 275546 600854
rect 275782 600618 275866 600854
rect 276102 600618 311546 600854
rect 311782 600618 311866 600854
rect 312102 600618 347546 600854
rect 347782 600618 347866 600854
rect 348102 600618 383546 600854
rect 383782 600618 383866 600854
rect 384102 600618 419546 600854
rect 419782 600618 419866 600854
rect 420102 600618 455546 600854
rect 455782 600618 455866 600854
rect 456102 600618 491546 600854
rect 491782 600618 491866 600854
rect 492102 600618 527546 600854
rect 527782 600618 527866 600854
rect 528102 600618 563546 600854
rect 563782 600618 563866 600854
rect 564102 600618 588222 600854
rect 588458 600618 588542 600854
rect 588778 600618 588810 600854
rect -4886 600586 588810 600618
rect -2966 597454 586890 597486
rect -2966 597218 -2934 597454
rect -2698 597218 -2614 597454
rect -2378 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 91826 597454
rect 92062 597218 92146 597454
rect 92382 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 163826 597454
rect 164062 597218 164146 597454
rect 164382 597218 199826 597454
rect 200062 597218 200146 597454
rect 200382 597218 235826 597454
rect 236062 597218 236146 597454
rect 236382 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 586302 597454
rect 586538 597218 586622 597454
rect 586858 597218 586890 597454
rect -2966 597134 586890 597218
rect -2966 596898 -2934 597134
rect -2698 596898 -2614 597134
rect -2378 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 91826 597134
rect 92062 596898 92146 597134
rect 92382 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 163826 597134
rect 164062 596898 164146 597134
rect 164382 596898 199826 597134
rect 200062 596898 200146 597134
rect 200382 596898 235826 597134
rect 236062 596898 236146 597134
rect 236382 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 586302 597134
rect 586538 596898 586622 597134
rect 586858 596898 586890 597134
rect -2966 596866 586890 596898
rect -8726 590614 592650 590646
rect -8726 590378 -7734 590614
rect -7498 590378 -7414 590614
rect -7178 590378 12986 590614
rect 13222 590378 13306 590614
rect 13542 590378 48986 590614
rect 49222 590378 49306 590614
rect 49542 590378 84986 590614
rect 85222 590378 85306 590614
rect 85542 590378 120986 590614
rect 121222 590378 121306 590614
rect 121542 590378 156986 590614
rect 157222 590378 157306 590614
rect 157542 590378 192986 590614
rect 193222 590378 193306 590614
rect 193542 590378 228986 590614
rect 229222 590378 229306 590614
rect 229542 590378 264986 590614
rect 265222 590378 265306 590614
rect 265542 590378 300986 590614
rect 301222 590378 301306 590614
rect 301542 590378 336986 590614
rect 337222 590378 337306 590614
rect 337542 590378 372986 590614
rect 373222 590378 373306 590614
rect 373542 590378 408986 590614
rect 409222 590378 409306 590614
rect 409542 590378 444986 590614
rect 445222 590378 445306 590614
rect 445542 590378 480986 590614
rect 481222 590378 481306 590614
rect 481542 590378 516986 590614
rect 517222 590378 517306 590614
rect 517542 590378 552986 590614
rect 553222 590378 553306 590614
rect 553542 590378 591102 590614
rect 591338 590378 591422 590614
rect 591658 590378 592650 590614
rect -8726 590294 592650 590378
rect -8726 590058 -7734 590294
rect -7498 590058 -7414 590294
rect -7178 590058 12986 590294
rect 13222 590058 13306 590294
rect 13542 590058 48986 590294
rect 49222 590058 49306 590294
rect 49542 590058 84986 590294
rect 85222 590058 85306 590294
rect 85542 590058 120986 590294
rect 121222 590058 121306 590294
rect 121542 590058 156986 590294
rect 157222 590058 157306 590294
rect 157542 590058 192986 590294
rect 193222 590058 193306 590294
rect 193542 590058 228986 590294
rect 229222 590058 229306 590294
rect 229542 590058 264986 590294
rect 265222 590058 265306 590294
rect 265542 590058 300986 590294
rect 301222 590058 301306 590294
rect 301542 590058 336986 590294
rect 337222 590058 337306 590294
rect 337542 590058 372986 590294
rect 373222 590058 373306 590294
rect 373542 590058 408986 590294
rect 409222 590058 409306 590294
rect 409542 590058 444986 590294
rect 445222 590058 445306 590294
rect 445542 590058 480986 590294
rect 481222 590058 481306 590294
rect 481542 590058 516986 590294
rect 517222 590058 517306 590294
rect 517542 590058 552986 590294
rect 553222 590058 553306 590294
rect 553542 590058 591102 590294
rect 591338 590058 591422 590294
rect 591658 590058 592650 590294
rect -8726 590026 592650 590058
rect -6806 586894 590730 586926
rect -6806 586658 -5814 586894
rect -5578 586658 -5494 586894
rect -5258 586658 9266 586894
rect 9502 586658 9586 586894
rect 9822 586658 45266 586894
rect 45502 586658 45586 586894
rect 45822 586658 81266 586894
rect 81502 586658 81586 586894
rect 81822 586658 117266 586894
rect 117502 586658 117586 586894
rect 117822 586658 153266 586894
rect 153502 586658 153586 586894
rect 153822 586658 189266 586894
rect 189502 586658 189586 586894
rect 189822 586658 225266 586894
rect 225502 586658 225586 586894
rect 225822 586658 261266 586894
rect 261502 586658 261586 586894
rect 261822 586658 297266 586894
rect 297502 586658 297586 586894
rect 297822 586658 333266 586894
rect 333502 586658 333586 586894
rect 333822 586658 369266 586894
rect 369502 586658 369586 586894
rect 369822 586658 405266 586894
rect 405502 586658 405586 586894
rect 405822 586658 441266 586894
rect 441502 586658 441586 586894
rect 441822 586658 477266 586894
rect 477502 586658 477586 586894
rect 477822 586658 513266 586894
rect 513502 586658 513586 586894
rect 513822 586658 549266 586894
rect 549502 586658 549586 586894
rect 549822 586658 589182 586894
rect 589418 586658 589502 586894
rect 589738 586658 590730 586894
rect -6806 586574 590730 586658
rect -6806 586338 -5814 586574
rect -5578 586338 -5494 586574
rect -5258 586338 9266 586574
rect 9502 586338 9586 586574
rect 9822 586338 45266 586574
rect 45502 586338 45586 586574
rect 45822 586338 81266 586574
rect 81502 586338 81586 586574
rect 81822 586338 117266 586574
rect 117502 586338 117586 586574
rect 117822 586338 153266 586574
rect 153502 586338 153586 586574
rect 153822 586338 189266 586574
rect 189502 586338 189586 586574
rect 189822 586338 225266 586574
rect 225502 586338 225586 586574
rect 225822 586338 261266 586574
rect 261502 586338 261586 586574
rect 261822 586338 297266 586574
rect 297502 586338 297586 586574
rect 297822 586338 333266 586574
rect 333502 586338 333586 586574
rect 333822 586338 369266 586574
rect 369502 586338 369586 586574
rect 369822 586338 405266 586574
rect 405502 586338 405586 586574
rect 405822 586338 441266 586574
rect 441502 586338 441586 586574
rect 441822 586338 477266 586574
rect 477502 586338 477586 586574
rect 477822 586338 513266 586574
rect 513502 586338 513586 586574
rect 513822 586338 549266 586574
rect 549502 586338 549586 586574
rect 549822 586338 589182 586574
rect 589418 586338 589502 586574
rect 589738 586338 590730 586574
rect -6806 586306 590730 586338
rect -4886 583174 588810 583206
rect -4886 582938 -3894 583174
rect -3658 582938 -3574 583174
rect -3338 582938 5546 583174
rect 5782 582938 5866 583174
rect 6102 582938 41546 583174
rect 41782 582938 41866 583174
rect 42102 582938 77546 583174
rect 77782 582938 77866 583174
rect 78102 582938 113546 583174
rect 113782 582938 113866 583174
rect 114102 582938 149546 583174
rect 149782 582938 149866 583174
rect 150102 582938 185546 583174
rect 185782 582938 185866 583174
rect 186102 582938 221546 583174
rect 221782 582938 221866 583174
rect 222102 582938 257546 583174
rect 257782 582938 257866 583174
rect 258102 582938 293546 583174
rect 293782 582938 293866 583174
rect 294102 582938 329546 583174
rect 329782 582938 329866 583174
rect 330102 582938 365546 583174
rect 365782 582938 365866 583174
rect 366102 582938 401546 583174
rect 401782 582938 401866 583174
rect 402102 582938 437546 583174
rect 437782 582938 437866 583174
rect 438102 582938 473546 583174
rect 473782 582938 473866 583174
rect 474102 582938 509546 583174
rect 509782 582938 509866 583174
rect 510102 582938 545546 583174
rect 545782 582938 545866 583174
rect 546102 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 587262 583174
rect 587498 582938 587582 583174
rect 587818 582938 588810 583174
rect -4886 582854 588810 582938
rect -4886 582618 -3894 582854
rect -3658 582618 -3574 582854
rect -3338 582618 5546 582854
rect 5782 582618 5866 582854
rect 6102 582618 41546 582854
rect 41782 582618 41866 582854
rect 42102 582618 77546 582854
rect 77782 582618 77866 582854
rect 78102 582618 113546 582854
rect 113782 582618 113866 582854
rect 114102 582618 149546 582854
rect 149782 582618 149866 582854
rect 150102 582618 185546 582854
rect 185782 582618 185866 582854
rect 186102 582618 221546 582854
rect 221782 582618 221866 582854
rect 222102 582618 257546 582854
rect 257782 582618 257866 582854
rect 258102 582618 293546 582854
rect 293782 582618 293866 582854
rect 294102 582618 329546 582854
rect 329782 582618 329866 582854
rect 330102 582618 365546 582854
rect 365782 582618 365866 582854
rect 366102 582618 401546 582854
rect 401782 582618 401866 582854
rect 402102 582618 437546 582854
rect 437782 582618 437866 582854
rect 438102 582618 473546 582854
rect 473782 582618 473866 582854
rect 474102 582618 509546 582854
rect 509782 582618 509866 582854
rect 510102 582618 545546 582854
rect 545782 582618 545866 582854
rect 546102 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 587262 582854
rect 587498 582618 587582 582854
rect 587818 582618 588810 582854
rect -4886 582586 588810 582618
rect -2966 579454 586890 579486
rect -2966 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 73826 579454
rect 74062 579218 74146 579454
rect 74382 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 586890 579454
rect -2966 579134 586890 579218
rect -2966 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 73826 579134
rect 74062 578898 74146 579134
rect 74382 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 586890 579134
rect -2966 578866 586890 578898
rect -8726 572614 592650 572646
rect -8726 572378 -8694 572614
rect -8458 572378 -8374 572614
rect -8138 572378 30986 572614
rect 31222 572378 31306 572614
rect 31542 572378 66986 572614
rect 67222 572378 67306 572614
rect 67542 572378 102986 572614
rect 103222 572378 103306 572614
rect 103542 572378 138986 572614
rect 139222 572378 139306 572614
rect 139542 572378 174986 572614
rect 175222 572378 175306 572614
rect 175542 572378 210986 572614
rect 211222 572378 211306 572614
rect 211542 572378 246986 572614
rect 247222 572378 247306 572614
rect 247542 572378 282986 572614
rect 283222 572378 283306 572614
rect 283542 572378 318986 572614
rect 319222 572378 319306 572614
rect 319542 572378 354986 572614
rect 355222 572378 355306 572614
rect 355542 572378 390986 572614
rect 391222 572378 391306 572614
rect 391542 572378 426986 572614
rect 427222 572378 427306 572614
rect 427542 572378 462986 572614
rect 463222 572378 463306 572614
rect 463542 572378 498986 572614
rect 499222 572378 499306 572614
rect 499542 572378 534986 572614
rect 535222 572378 535306 572614
rect 535542 572378 570986 572614
rect 571222 572378 571306 572614
rect 571542 572378 592062 572614
rect 592298 572378 592382 572614
rect 592618 572378 592650 572614
rect -8726 572294 592650 572378
rect -8726 572058 -8694 572294
rect -8458 572058 -8374 572294
rect -8138 572058 30986 572294
rect 31222 572058 31306 572294
rect 31542 572058 66986 572294
rect 67222 572058 67306 572294
rect 67542 572058 102986 572294
rect 103222 572058 103306 572294
rect 103542 572058 138986 572294
rect 139222 572058 139306 572294
rect 139542 572058 174986 572294
rect 175222 572058 175306 572294
rect 175542 572058 210986 572294
rect 211222 572058 211306 572294
rect 211542 572058 246986 572294
rect 247222 572058 247306 572294
rect 247542 572058 282986 572294
rect 283222 572058 283306 572294
rect 283542 572058 318986 572294
rect 319222 572058 319306 572294
rect 319542 572058 354986 572294
rect 355222 572058 355306 572294
rect 355542 572058 390986 572294
rect 391222 572058 391306 572294
rect 391542 572058 426986 572294
rect 427222 572058 427306 572294
rect 427542 572058 462986 572294
rect 463222 572058 463306 572294
rect 463542 572058 498986 572294
rect 499222 572058 499306 572294
rect 499542 572058 534986 572294
rect 535222 572058 535306 572294
rect 535542 572058 570986 572294
rect 571222 572058 571306 572294
rect 571542 572058 592062 572294
rect 592298 572058 592382 572294
rect 592618 572058 592650 572294
rect -8726 572026 592650 572058
rect -6806 568894 590730 568926
rect -6806 568658 -6774 568894
rect -6538 568658 -6454 568894
rect -6218 568658 27266 568894
rect 27502 568658 27586 568894
rect 27822 568658 63266 568894
rect 63502 568658 63586 568894
rect 63822 568658 99266 568894
rect 99502 568658 99586 568894
rect 99822 568658 135266 568894
rect 135502 568658 135586 568894
rect 135822 568658 171266 568894
rect 171502 568658 171586 568894
rect 171822 568658 207266 568894
rect 207502 568658 207586 568894
rect 207822 568658 243266 568894
rect 243502 568658 243586 568894
rect 243822 568658 279266 568894
rect 279502 568658 279586 568894
rect 279822 568658 315266 568894
rect 315502 568658 315586 568894
rect 315822 568658 351266 568894
rect 351502 568658 351586 568894
rect 351822 568658 387266 568894
rect 387502 568658 387586 568894
rect 387822 568658 423266 568894
rect 423502 568658 423586 568894
rect 423822 568658 459266 568894
rect 459502 568658 459586 568894
rect 459822 568658 495266 568894
rect 495502 568658 495586 568894
rect 495822 568658 531266 568894
rect 531502 568658 531586 568894
rect 531822 568658 567266 568894
rect 567502 568658 567586 568894
rect 567822 568658 590142 568894
rect 590378 568658 590462 568894
rect 590698 568658 590730 568894
rect -6806 568574 590730 568658
rect -6806 568338 -6774 568574
rect -6538 568338 -6454 568574
rect -6218 568338 27266 568574
rect 27502 568338 27586 568574
rect 27822 568338 63266 568574
rect 63502 568338 63586 568574
rect 63822 568338 99266 568574
rect 99502 568338 99586 568574
rect 99822 568338 135266 568574
rect 135502 568338 135586 568574
rect 135822 568338 171266 568574
rect 171502 568338 171586 568574
rect 171822 568338 207266 568574
rect 207502 568338 207586 568574
rect 207822 568338 243266 568574
rect 243502 568338 243586 568574
rect 243822 568338 279266 568574
rect 279502 568338 279586 568574
rect 279822 568338 315266 568574
rect 315502 568338 315586 568574
rect 315822 568338 351266 568574
rect 351502 568338 351586 568574
rect 351822 568338 387266 568574
rect 387502 568338 387586 568574
rect 387822 568338 423266 568574
rect 423502 568338 423586 568574
rect 423822 568338 459266 568574
rect 459502 568338 459586 568574
rect 459822 568338 495266 568574
rect 495502 568338 495586 568574
rect 495822 568338 531266 568574
rect 531502 568338 531586 568574
rect 531822 568338 567266 568574
rect 567502 568338 567586 568574
rect 567822 568338 590142 568574
rect 590378 568338 590462 568574
rect 590698 568338 590730 568574
rect -6806 568306 590730 568338
rect -4886 565174 588810 565206
rect -4886 564938 -4854 565174
rect -4618 564938 -4534 565174
rect -4298 564938 23546 565174
rect 23782 564938 23866 565174
rect 24102 564938 59546 565174
rect 59782 564938 59866 565174
rect 60102 564938 95546 565174
rect 95782 564938 95866 565174
rect 96102 564938 131546 565174
rect 131782 564938 131866 565174
rect 132102 564938 167546 565174
rect 167782 564938 167866 565174
rect 168102 564938 203546 565174
rect 203782 564938 203866 565174
rect 204102 564938 239546 565174
rect 239782 564938 239866 565174
rect 240102 564938 275546 565174
rect 275782 564938 275866 565174
rect 276102 564938 311546 565174
rect 311782 564938 311866 565174
rect 312102 564938 347546 565174
rect 347782 564938 347866 565174
rect 348102 564938 383546 565174
rect 383782 564938 383866 565174
rect 384102 564938 419546 565174
rect 419782 564938 419866 565174
rect 420102 564938 455546 565174
rect 455782 564938 455866 565174
rect 456102 564938 491546 565174
rect 491782 564938 491866 565174
rect 492102 564938 527546 565174
rect 527782 564938 527866 565174
rect 528102 564938 563546 565174
rect 563782 564938 563866 565174
rect 564102 564938 588222 565174
rect 588458 564938 588542 565174
rect 588778 564938 588810 565174
rect -4886 564854 588810 564938
rect -4886 564618 -4854 564854
rect -4618 564618 -4534 564854
rect -4298 564618 23546 564854
rect 23782 564618 23866 564854
rect 24102 564618 59546 564854
rect 59782 564618 59866 564854
rect 60102 564618 95546 564854
rect 95782 564618 95866 564854
rect 96102 564618 131546 564854
rect 131782 564618 131866 564854
rect 132102 564618 167546 564854
rect 167782 564618 167866 564854
rect 168102 564618 203546 564854
rect 203782 564618 203866 564854
rect 204102 564618 239546 564854
rect 239782 564618 239866 564854
rect 240102 564618 275546 564854
rect 275782 564618 275866 564854
rect 276102 564618 311546 564854
rect 311782 564618 311866 564854
rect 312102 564618 347546 564854
rect 347782 564618 347866 564854
rect 348102 564618 383546 564854
rect 383782 564618 383866 564854
rect 384102 564618 419546 564854
rect 419782 564618 419866 564854
rect 420102 564618 455546 564854
rect 455782 564618 455866 564854
rect 456102 564618 491546 564854
rect 491782 564618 491866 564854
rect 492102 564618 527546 564854
rect 527782 564618 527866 564854
rect 528102 564618 563546 564854
rect 563782 564618 563866 564854
rect 564102 564618 588222 564854
rect 588458 564618 588542 564854
rect 588778 564618 588810 564854
rect -4886 564586 588810 564618
rect -2966 561454 586890 561486
rect -2966 561218 -2934 561454
rect -2698 561218 -2614 561454
rect -2378 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 91826 561454
rect 92062 561218 92146 561454
rect 92382 561218 127826 561454
rect 128062 561218 128146 561454
rect 128382 561218 163826 561454
rect 164062 561218 164146 561454
rect 164382 561218 199826 561454
rect 200062 561218 200146 561454
rect 200382 561218 235826 561454
rect 236062 561218 236146 561454
rect 236382 561218 271826 561454
rect 272062 561218 272146 561454
rect 272382 561218 307826 561454
rect 308062 561218 308146 561454
rect 308382 561218 343826 561454
rect 344062 561218 344146 561454
rect 344382 561218 379826 561454
rect 380062 561218 380146 561454
rect 380382 561218 415826 561454
rect 416062 561218 416146 561454
rect 416382 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 586302 561454
rect 586538 561218 586622 561454
rect 586858 561218 586890 561454
rect -2966 561134 586890 561218
rect -2966 560898 -2934 561134
rect -2698 560898 -2614 561134
rect -2378 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 91826 561134
rect 92062 560898 92146 561134
rect 92382 560898 127826 561134
rect 128062 560898 128146 561134
rect 128382 560898 163826 561134
rect 164062 560898 164146 561134
rect 164382 560898 199826 561134
rect 200062 560898 200146 561134
rect 200382 560898 235826 561134
rect 236062 560898 236146 561134
rect 236382 560898 271826 561134
rect 272062 560898 272146 561134
rect 272382 560898 307826 561134
rect 308062 560898 308146 561134
rect 308382 560898 343826 561134
rect 344062 560898 344146 561134
rect 344382 560898 379826 561134
rect 380062 560898 380146 561134
rect 380382 560898 415826 561134
rect 416062 560898 416146 561134
rect 416382 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 586302 561134
rect 586538 560898 586622 561134
rect 586858 560898 586890 561134
rect -2966 560866 586890 560898
rect -8726 554614 592650 554646
rect -8726 554378 -7734 554614
rect -7498 554378 -7414 554614
rect -7178 554378 12986 554614
rect 13222 554378 13306 554614
rect 13542 554378 48986 554614
rect 49222 554378 49306 554614
rect 49542 554378 84986 554614
rect 85222 554378 85306 554614
rect 85542 554378 120986 554614
rect 121222 554378 121306 554614
rect 121542 554378 156986 554614
rect 157222 554378 157306 554614
rect 157542 554378 192986 554614
rect 193222 554378 193306 554614
rect 193542 554378 228986 554614
rect 229222 554378 229306 554614
rect 229542 554378 264986 554614
rect 265222 554378 265306 554614
rect 265542 554378 300986 554614
rect 301222 554378 301306 554614
rect 301542 554378 336986 554614
rect 337222 554378 337306 554614
rect 337542 554378 372986 554614
rect 373222 554378 373306 554614
rect 373542 554378 408986 554614
rect 409222 554378 409306 554614
rect 409542 554378 444986 554614
rect 445222 554378 445306 554614
rect 445542 554378 480986 554614
rect 481222 554378 481306 554614
rect 481542 554378 516986 554614
rect 517222 554378 517306 554614
rect 517542 554378 552986 554614
rect 553222 554378 553306 554614
rect 553542 554378 591102 554614
rect 591338 554378 591422 554614
rect 591658 554378 592650 554614
rect -8726 554294 592650 554378
rect -8726 554058 -7734 554294
rect -7498 554058 -7414 554294
rect -7178 554058 12986 554294
rect 13222 554058 13306 554294
rect 13542 554058 48986 554294
rect 49222 554058 49306 554294
rect 49542 554058 84986 554294
rect 85222 554058 85306 554294
rect 85542 554058 120986 554294
rect 121222 554058 121306 554294
rect 121542 554058 156986 554294
rect 157222 554058 157306 554294
rect 157542 554058 192986 554294
rect 193222 554058 193306 554294
rect 193542 554058 228986 554294
rect 229222 554058 229306 554294
rect 229542 554058 264986 554294
rect 265222 554058 265306 554294
rect 265542 554058 300986 554294
rect 301222 554058 301306 554294
rect 301542 554058 336986 554294
rect 337222 554058 337306 554294
rect 337542 554058 372986 554294
rect 373222 554058 373306 554294
rect 373542 554058 408986 554294
rect 409222 554058 409306 554294
rect 409542 554058 444986 554294
rect 445222 554058 445306 554294
rect 445542 554058 480986 554294
rect 481222 554058 481306 554294
rect 481542 554058 516986 554294
rect 517222 554058 517306 554294
rect 517542 554058 552986 554294
rect 553222 554058 553306 554294
rect 553542 554058 591102 554294
rect 591338 554058 591422 554294
rect 591658 554058 592650 554294
rect -8726 554026 592650 554058
rect -6806 550894 590730 550926
rect -6806 550658 -5814 550894
rect -5578 550658 -5494 550894
rect -5258 550658 9266 550894
rect 9502 550658 9586 550894
rect 9822 550658 45266 550894
rect 45502 550658 45586 550894
rect 45822 550658 81266 550894
rect 81502 550658 81586 550894
rect 81822 550658 117266 550894
rect 117502 550658 117586 550894
rect 117822 550658 153266 550894
rect 153502 550658 153586 550894
rect 153822 550658 189266 550894
rect 189502 550658 189586 550894
rect 189822 550658 225266 550894
rect 225502 550658 225586 550894
rect 225822 550658 261266 550894
rect 261502 550658 261586 550894
rect 261822 550658 297266 550894
rect 297502 550658 297586 550894
rect 297822 550658 333266 550894
rect 333502 550658 333586 550894
rect 333822 550658 369266 550894
rect 369502 550658 369586 550894
rect 369822 550658 405266 550894
rect 405502 550658 405586 550894
rect 405822 550658 441266 550894
rect 441502 550658 441586 550894
rect 441822 550658 477266 550894
rect 477502 550658 477586 550894
rect 477822 550658 513266 550894
rect 513502 550658 513586 550894
rect 513822 550658 549266 550894
rect 549502 550658 549586 550894
rect 549822 550658 589182 550894
rect 589418 550658 589502 550894
rect 589738 550658 590730 550894
rect -6806 550574 590730 550658
rect -6806 550338 -5814 550574
rect -5578 550338 -5494 550574
rect -5258 550338 9266 550574
rect 9502 550338 9586 550574
rect 9822 550338 45266 550574
rect 45502 550338 45586 550574
rect 45822 550338 81266 550574
rect 81502 550338 81586 550574
rect 81822 550338 117266 550574
rect 117502 550338 117586 550574
rect 117822 550338 153266 550574
rect 153502 550338 153586 550574
rect 153822 550338 189266 550574
rect 189502 550338 189586 550574
rect 189822 550338 225266 550574
rect 225502 550338 225586 550574
rect 225822 550338 261266 550574
rect 261502 550338 261586 550574
rect 261822 550338 297266 550574
rect 297502 550338 297586 550574
rect 297822 550338 333266 550574
rect 333502 550338 333586 550574
rect 333822 550338 369266 550574
rect 369502 550338 369586 550574
rect 369822 550338 405266 550574
rect 405502 550338 405586 550574
rect 405822 550338 441266 550574
rect 441502 550338 441586 550574
rect 441822 550338 477266 550574
rect 477502 550338 477586 550574
rect 477822 550338 513266 550574
rect 513502 550338 513586 550574
rect 513822 550338 549266 550574
rect 549502 550338 549586 550574
rect 549822 550338 589182 550574
rect 589418 550338 589502 550574
rect 589738 550338 590730 550574
rect -6806 550306 590730 550338
rect -4886 547174 588810 547206
rect -4886 546938 -3894 547174
rect -3658 546938 -3574 547174
rect -3338 546938 5546 547174
rect 5782 546938 5866 547174
rect 6102 546938 41546 547174
rect 41782 546938 41866 547174
rect 42102 546938 77546 547174
rect 77782 546938 77866 547174
rect 78102 546938 113546 547174
rect 113782 546938 113866 547174
rect 114102 546938 149546 547174
rect 149782 546938 149866 547174
rect 150102 546938 185546 547174
rect 185782 546938 185866 547174
rect 186102 546938 221546 547174
rect 221782 546938 221866 547174
rect 222102 546938 257546 547174
rect 257782 546938 257866 547174
rect 258102 546938 293546 547174
rect 293782 546938 293866 547174
rect 294102 546938 329546 547174
rect 329782 546938 329866 547174
rect 330102 546938 365546 547174
rect 365782 546938 365866 547174
rect 366102 546938 401546 547174
rect 401782 546938 401866 547174
rect 402102 546938 437546 547174
rect 437782 546938 437866 547174
rect 438102 546938 473546 547174
rect 473782 546938 473866 547174
rect 474102 546938 509546 547174
rect 509782 546938 509866 547174
rect 510102 546938 545546 547174
rect 545782 546938 545866 547174
rect 546102 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 587262 547174
rect 587498 546938 587582 547174
rect 587818 546938 588810 547174
rect -4886 546854 588810 546938
rect -4886 546618 -3894 546854
rect -3658 546618 -3574 546854
rect -3338 546618 5546 546854
rect 5782 546618 5866 546854
rect 6102 546618 41546 546854
rect 41782 546618 41866 546854
rect 42102 546618 77546 546854
rect 77782 546618 77866 546854
rect 78102 546618 113546 546854
rect 113782 546618 113866 546854
rect 114102 546618 149546 546854
rect 149782 546618 149866 546854
rect 150102 546618 185546 546854
rect 185782 546618 185866 546854
rect 186102 546618 221546 546854
rect 221782 546618 221866 546854
rect 222102 546618 257546 546854
rect 257782 546618 257866 546854
rect 258102 546618 293546 546854
rect 293782 546618 293866 546854
rect 294102 546618 329546 546854
rect 329782 546618 329866 546854
rect 330102 546618 365546 546854
rect 365782 546618 365866 546854
rect 366102 546618 401546 546854
rect 401782 546618 401866 546854
rect 402102 546618 437546 546854
rect 437782 546618 437866 546854
rect 438102 546618 473546 546854
rect 473782 546618 473866 546854
rect 474102 546618 509546 546854
rect 509782 546618 509866 546854
rect 510102 546618 545546 546854
rect 545782 546618 545866 546854
rect 546102 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 587262 546854
rect 587498 546618 587582 546854
rect 587818 546618 588810 546854
rect -4886 546586 588810 546618
rect -2966 543454 586890 543486
rect -2966 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 73826 543454
rect 74062 543218 74146 543454
rect 74382 543218 109826 543454
rect 110062 543218 110146 543454
rect 110382 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 217826 543454
rect 218062 543218 218146 543454
rect 218382 543218 253826 543454
rect 254062 543218 254146 543454
rect 254382 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 325826 543454
rect 326062 543218 326146 543454
rect 326382 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 586890 543454
rect -2966 543134 586890 543218
rect -2966 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 73826 543134
rect 74062 542898 74146 543134
rect 74382 542898 109826 543134
rect 110062 542898 110146 543134
rect 110382 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 217826 543134
rect 218062 542898 218146 543134
rect 218382 542898 253826 543134
rect 254062 542898 254146 543134
rect 254382 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 325826 543134
rect 326062 542898 326146 543134
rect 326382 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 586890 543134
rect -2966 542866 586890 542898
rect -8726 536614 592650 536646
rect -8726 536378 -8694 536614
rect -8458 536378 -8374 536614
rect -8138 536378 30986 536614
rect 31222 536378 31306 536614
rect 31542 536378 66986 536614
rect 67222 536378 67306 536614
rect 67542 536378 102986 536614
rect 103222 536378 103306 536614
rect 103542 536378 138986 536614
rect 139222 536378 139306 536614
rect 139542 536378 174986 536614
rect 175222 536378 175306 536614
rect 175542 536378 210986 536614
rect 211222 536378 211306 536614
rect 211542 536378 246986 536614
rect 247222 536378 247306 536614
rect 247542 536378 282986 536614
rect 283222 536378 283306 536614
rect 283542 536378 318986 536614
rect 319222 536378 319306 536614
rect 319542 536378 354986 536614
rect 355222 536378 355306 536614
rect 355542 536378 390986 536614
rect 391222 536378 391306 536614
rect 391542 536378 426986 536614
rect 427222 536378 427306 536614
rect 427542 536378 462986 536614
rect 463222 536378 463306 536614
rect 463542 536378 498986 536614
rect 499222 536378 499306 536614
rect 499542 536378 534986 536614
rect 535222 536378 535306 536614
rect 535542 536378 570986 536614
rect 571222 536378 571306 536614
rect 571542 536378 592062 536614
rect 592298 536378 592382 536614
rect 592618 536378 592650 536614
rect -8726 536294 592650 536378
rect -8726 536058 -8694 536294
rect -8458 536058 -8374 536294
rect -8138 536058 30986 536294
rect 31222 536058 31306 536294
rect 31542 536058 66986 536294
rect 67222 536058 67306 536294
rect 67542 536058 102986 536294
rect 103222 536058 103306 536294
rect 103542 536058 138986 536294
rect 139222 536058 139306 536294
rect 139542 536058 174986 536294
rect 175222 536058 175306 536294
rect 175542 536058 210986 536294
rect 211222 536058 211306 536294
rect 211542 536058 246986 536294
rect 247222 536058 247306 536294
rect 247542 536058 282986 536294
rect 283222 536058 283306 536294
rect 283542 536058 318986 536294
rect 319222 536058 319306 536294
rect 319542 536058 354986 536294
rect 355222 536058 355306 536294
rect 355542 536058 390986 536294
rect 391222 536058 391306 536294
rect 391542 536058 426986 536294
rect 427222 536058 427306 536294
rect 427542 536058 462986 536294
rect 463222 536058 463306 536294
rect 463542 536058 498986 536294
rect 499222 536058 499306 536294
rect 499542 536058 534986 536294
rect 535222 536058 535306 536294
rect 535542 536058 570986 536294
rect 571222 536058 571306 536294
rect 571542 536058 592062 536294
rect 592298 536058 592382 536294
rect 592618 536058 592650 536294
rect -8726 536026 592650 536058
rect -6806 532894 590730 532926
rect -6806 532658 -6774 532894
rect -6538 532658 -6454 532894
rect -6218 532658 27266 532894
rect 27502 532658 27586 532894
rect 27822 532658 63266 532894
rect 63502 532658 63586 532894
rect 63822 532658 99266 532894
rect 99502 532658 99586 532894
rect 99822 532658 135266 532894
rect 135502 532658 135586 532894
rect 135822 532658 171266 532894
rect 171502 532658 171586 532894
rect 171822 532658 207266 532894
rect 207502 532658 207586 532894
rect 207822 532658 243266 532894
rect 243502 532658 243586 532894
rect 243822 532658 279266 532894
rect 279502 532658 279586 532894
rect 279822 532658 315266 532894
rect 315502 532658 315586 532894
rect 315822 532658 351266 532894
rect 351502 532658 351586 532894
rect 351822 532658 387266 532894
rect 387502 532658 387586 532894
rect 387822 532658 423266 532894
rect 423502 532658 423586 532894
rect 423822 532658 459266 532894
rect 459502 532658 459586 532894
rect 459822 532658 495266 532894
rect 495502 532658 495586 532894
rect 495822 532658 531266 532894
rect 531502 532658 531586 532894
rect 531822 532658 567266 532894
rect 567502 532658 567586 532894
rect 567822 532658 590142 532894
rect 590378 532658 590462 532894
rect 590698 532658 590730 532894
rect -6806 532574 590730 532658
rect -6806 532338 -6774 532574
rect -6538 532338 -6454 532574
rect -6218 532338 27266 532574
rect 27502 532338 27586 532574
rect 27822 532338 63266 532574
rect 63502 532338 63586 532574
rect 63822 532338 99266 532574
rect 99502 532338 99586 532574
rect 99822 532338 135266 532574
rect 135502 532338 135586 532574
rect 135822 532338 171266 532574
rect 171502 532338 171586 532574
rect 171822 532338 207266 532574
rect 207502 532338 207586 532574
rect 207822 532338 243266 532574
rect 243502 532338 243586 532574
rect 243822 532338 279266 532574
rect 279502 532338 279586 532574
rect 279822 532338 315266 532574
rect 315502 532338 315586 532574
rect 315822 532338 351266 532574
rect 351502 532338 351586 532574
rect 351822 532338 387266 532574
rect 387502 532338 387586 532574
rect 387822 532338 423266 532574
rect 423502 532338 423586 532574
rect 423822 532338 459266 532574
rect 459502 532338 459586 532574
rect 459822 532338 495266 532574
rect 495502 532338 495586 532574
rect 495822 532338 531266 532574
rect 531502 532338 531586 532574
rect 531822 532338 567266 532574
rect 567502 532338 567586 532574
rect 567822 532338 590142 532574
rect 590378 532338 590462 532574
rect 590698 532338 590730 532574
rect -6806 532306 590730 532338
rect -4886 529174 588810 529206
rect -4886 528938 -4854 529174
rect -4618 528938 -4534 529174
rect -4298 528938 23546 529174
rect 23782 528938 23866 529174
rect 24102 528938 59546 529174
rect 59782 528938 59866 529174
rect 60102 528938 95546 529174
rect 95782 528938 95866 529174
rect 96102 528938 131546 529174
rect 131782 528938 131866 529174
rect 132102 528938 167546 529174
rect 167782 528938 167866 529174
rect 168102 528938 203546 529174
rect 203782 528938 203866 529174
rect 204102 528938 239546 529174
rect 239782 528938 239866 529174
rect 240102 528938 275546 529174
rect 275782 528938 275866 529174
rect 276102 528938 311546 529174
rect 311782 528938 311866 529174
rect 312102 528938 347546 529174
rect 347782 528938 347866 529174
rect 348102 528938 383546 529174
rect 383782 528938 383866 529174
rect 384102 528938 419546 529174
rect 419782 528938 419866 529174
rect 420102 528938 455546 529174
rect 455782 528938 455866 529174
rect 456102 528938 491546 529174
rect 491782 528938 491866 529174
rect 492102 528938 527546 529174
rect 527782 528938 527866 529174
rect 528102 528938 563546 529174
rect 563782 528938 563866 529174
rect 564102 528938 588222 529174
rect 588458 528938 588542 529174
rect 588778 528938 588810 529174
rect -4886 528854 588810 528938
rect -4886 528618 -4854 528854
rect -4618 528618 -4534 528854
rect -4298 528618 23546 528854
rect 23782 528618 23866 528854
rect 24102 528618 59546 528854
rect 59782 528618 59866 528854
rect 60102 528618 95546 528854
rect 95782 528618 95866 528854
rect 96102 528618 131546 528854
rect 131782 528618 131866 528854
rect 132102 528618 167546 528854
rect 167782 528618 167866 528854
rect 168102 528618 203546 528854
rect 203782 528618 203866 528854
rect 204102 528618 239546 528854
rect 239782 528618 239866 528854
rect 240102 528618 275546 528854
rect 275782 528618 275866 528854
rect 276102 528618 311546 528854
rect 311782 528618 311866 528854
rect 312102 528618 347546 528854
rect 347782 528618 347866 528854
rect 348102 528618 383546 528854
rect 383782 528618 383866 528854
rect 384102 528618 419546 528854
rect 419782 528618 419866 528854
rect 420102 528618 455546 528854
rect 455782 528618 455866 528854
rect 456102 528618 491546 528854
rect 491782 528618 491866 528854
rect 492102 528618 527546 528854
rect 527782 528618 527866 528854
rect 528102 528618 563546 528854
rect 563782 528618 563866 528854
rect 564102 528618 588222 528854
rect 588458 528618 588542 528854
rect 588778 528618 588810 528854
rect -4886 528586 588810 528618
rect -2966 525454 586890 525486
rect -2966 525218 -2934 525454
rect -2698 525218 -2614 525454
rect -2378 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 91826 525454
rect 92062 525218 92146 525454
rect 92382 525218 127826 525454
rect 128062 525218 128146 525454
rect 128382 525218 163826 525454
rect 164062 525218 164146 525454
rect 164382 525218 199826 525454
rect 200062 525218 200146 525454
rect 200382 525218 235826 525454
rect 236062 525218 236146 525454
rect 236382 525218 271826 525454
rect 272062 525218 272146 525454
rect 272382 525218 307826 525454
rect 308062 525218 308146 525454
rect 308382 525218 343826 525454
rect 344062 525218 344146 525454
rect 344382 525218 379826 525454
rect 380062 525218 380146 525454
rect 380382 525218 415826 525454
rect 416062 525218 416146 525454
rect 416382 525218 451826 525454
rect 452062 525218 452146 525454
rect 452382 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 586302 525454
rect 586538 525218 586622 525454
rect 586858 525218 586890 525454
rect -2966 525134 586890 525218
rect -2966 524898 -2934 525134
rect -2698 524898 -2614 525134
rect -2378 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 91826 525134
rect 92062 524898 92146 525134
rect 92382 524898 127826 525134
rect 128062 524898 128146 525134
rect 128382 524898 163826 525134
rect 164062 524898 164146 525134
rect 164382 524898 199826 525134
rect 200062 524898 200146 525134
rect 200382 524898 235826 525134
rect 236062 524898 236146 525134
rect 236382 524898 271826 525134
rect 272062 524898 272146 525134
rect 272382 524898 307826 525134
rect 308062 524898 308146 525134
rect 308382 524898 343826 525134
rect 344062 524898 344146 525134
rect 344382 524898 379826 525134
rect 380062 524898 380146 525134
rect 380382 524898 415826 525134
rect 416062 524898 416146 525134
rect 416382 524898 451826 525134
rect 452062 524898 452146 525134
rect 452382 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 586302 525134
rect 586538 524898 586622 525134
rect 586858 524898 586890 525134
rect -2966 524866 586890 524898
rect -8726 518614 592650 518646
rect -8726 518378 -7734 518614
rect -7498 518378 -7414 518614
rect -7178 518378 12986 518614
rect 13222 518378 13306 518614
rect 13542 518378 48986 518614
rect 49222 518378 49306 518614
rect 49542 518378 84986 518614
rect 85222 518378 85306 518614
rect 85542 518378 120986 518614
rect 121222 518378 121306 518614
rect 121542 518378 156986 518614
rect 157222 518378 157306 518614
rect 157542 518378 192986 518614
rect 193222 518378 193306 518614
rect 193542 518378 228986 518614
rect 229222 518378 229306 518614
rect 229542 518378 264986 518614
rect 265222 518378 265306 518614
rect 265542 518378 300986 518614
rect 301222 518378 301306 518614
rect 301542 518378 336986 518614
rect 337222 518378 337306 518614
rect 337542 518378 372986 518614
rect 373222 518378 373306 518614
rect 373542 518378 408986 518614
rect 409222 518378 409306 518614
rect 409542 518378 444986 518614
rect 445222 518378 445306 518614
rect 445542 518378 480986 518614
rect 481222 518378 481306 518614
rect 481542 518378 516986 518614
rect 517222 518378 517306 518614
rect 517542 518378 552986 518614
rect 553222 518378 553306 518614
rect 553542 518378 591102 518614
rect 591338 518378 591422 518614
rect 591658 518378 592650 518614
rect -8726 518294 592650 518378
rect -8726 518058 -7734 518294
rect -7498 518058 -7414 518294
rect -7178 518058 12986 518294
rect 13222 518058 13306 518294
rect 13542 518058 48986 518294
rect 49222 518058 49306 518294
rect 49542 518058 84986 518294
rect 85222 518058 85306 518294
rect 85542 518058 120986 518294
rect 121222 518058 121306 518294
rect 121542 518058 156986 518294
rect 157222 518058 157306 518294
rect 157542 518058 192986 518294
rect 193222 518058 193306 518294
rect 193542 518058 228986 518294
rect 229222 518058 229306 518294
rect 229542 518058 264986 518294
rect 265222 518058 265306 518294
rect 265542 518058 300986 518294
rect 301222 518058 301306 518294
rect 301542 518058 336986 518294
rect 337222 518058 337306 518294
rect 337542 518058 372986 518294
rect 373222 518058 373306 518294
rect 373542 518058 408986 518294
rect 409222 518058 409306 518294
rect 409542 518058 444986 518294
rect 445222 518058 445306 518294
rect 445542 518058 480986 518294
rect 481222 518058 481306 518294
rect 481542 518058 516986 518294
rect 517222 518058 517306 518294
rect 517542 518058 552986 518294
rect 553222 518058 553306 518294
rect 553542 518058 591102 518294
rect 591338 518058 591422 518294
rect 591658 518058 592650 518294
rect -8726 518026 592650 518058
rect -6806 514894 590730 514926
rect -6806 514658 -5814 514894
rect -5578 514658 -5494 514894
rect -5258 514658 9266 514894
rect 9502 514658 9586 514894
rect 9822 514658 45266 514894
rect 45502 514658 45586 514894
rect 45822 514658 81266 514894
rect 81502 514658 81586 514894
rect 81822 514658 117266 514894
rect 117502 514658 117586 514894
rect 117822 514658 153266 514894
rect 153502 514658 153586 514894
rect 153822 514658 189266 514894
rect 189502 514658 189586 514894
rect 189822 514658 225266 514894
rect 225502 514658 225586 514894
rect 225822 514658 261266 514894
rect 261502 514658 261586 514894
rect 261822 514658 297266 514894
rect 297502 514658 297586 514894
rect 297822 514658 333266 514894
rect 333502 514658 333586 514894
rect 333822 514658 369266 514894
rect 369502 514658 369586 514894
rect 369822 514658 405266 514894
rect 405502 514658 405586 514894
rect 405822 514658 441266 514894
rect 441502 514658 441586 514894
rect 441822 514658 477266 514894
rect 477502 514658 477586 514894
rect 477822 514658 513266 514894
rect 513502 514658 513586 514894
rect 513822 514658 549266 514894
rect 549502 514658 549586 514894
rect 549822 514658 589182 514894
rect 589418 514658 589502 514894
rect 589738 514658 590730 514894
rect -6806 514574 590730 514658
rect -6806 514338 -5814 514574
rect -5578 514338 -5494 514574
rect -5258 514338 9266 514574
rect 9502 514338 9586 514574
rect 9822 514338 45266 514574
rect 45502 514338 45586 514574
rect 45822 514338 81266 514574
rect 81502 514338 81586 514574
rect 81822 514338 117266 514574
rect 117502 514338 117586 514574
rect 117822 514338 153266 514574
rect 153502 514338 153586 514574
rect 153822 514338 189266 514574
rect 189502 514338 189586 514574
rect 189822 514338 225266 514574
rect 225502 514338 225586 514574
rect 225822 514338 261266 514574
rect 261502 514338 261586 514574
rect 261822 514338 297266 514574
rect 297502 514338 297586 514574
rect 297822 514338 333266 514574
rect 333502 514338 333586 514574
rect 333822 514338 369266 514574
rect 369502 514338 369586 514574
rect 369822 514338 405266 514574
rect 405502 514338 405586 514574
rect 405822 514338 441266 514574
rect 441502 514338 441586 514574
rect 441822 514338 477266 514574
rect 477502 514338 477586 514574
rect 477822 514338 513266 514574
rect 513502 514338 513586 514574
rect 513822 514338 549266 514574
rect 549502 514338 549586 514574
rect 549822 514338 589182 514574
rect 589418 514338 589502 514574
rect 589738 514338 590730 514574
rect -6806 514306 590730 514338
rect -4886 511174 588810 511206
rect -4886 510938 -3894 511174
rect -3658 510938 -3574 511174
rect -3338 510938 5546 511174
rect 5782 510938 5866 511174
rect 6102 510938 41546 511174
rect 41782 510938 41866 511174
rect 42102 510938 77546 511174
rect 77782 510938 77866 511174
rect 78102 510938 113546 511174
rect 113782 510938 113866 511174
rect 114102 510938 149546 511174
rect 149782 510938 149866 511174
rect 150102 510938 185546 511174
rect 185782 510938 185866 511174
rect 186102 510938 221546 511174
rect 221782 510938 221866 511174
rect 222102 510938 257546 511174
rect 257782 510938 257866 511174
rect 258102 510938 293546 511174
rect 293782 510938 293866 511174
rect 294102 510938 329546 511174
rect 329782 510938 329866 511174
rect 330102 510938 365546 511174
rect 365782 510938 365866 511174
rect 366102 510938 401546 511174
rect 401782 510938 401866 511174
rect 402102 510938 437546 511174
rect 437782 510938 437866 511174
rect 438102 510938 473546 511174
rect 473782 510938 473866 511174
rect 474102 510938 509546 511174
rect 509782 510938 509866 511174
rect 510102 510938 545546 511174
rect 545782 510938 545866 511174
rect 546102 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 587262 511174
rect 587498 510938 587582 511174
rect 587818 510938 588810 511174
rect -4886 510854 588810 510938
rect -4886 510618 -3894 510854
rect -3658 510618 -3574 510854
rect -3338 510618 5546 510854
rect 5782 510618 5866 510854
rect 6102 510618 41546 510854
rect 41782 510618 41866 510854
rect 42102 510618 77546 510854
rect 77782 510618 77866 510854
rect 78102 510618 113546 510854
rect 113782 510618 113866 510854
rect 114102 510618 149546 510854
rect 149782 510618 149866 510854
rect 150102 510618 185546 510854
rect 185782 510618 185866 510854
rect 186102 510618 221546 510854
rect 221782 510618 221866 510854
rect 222102 510618 257546 510854
rect 257782 510618 257866 510854
rect 258102 510618 293546 510854
rect 293782 510618 293866 510854
rect 294102 510618 329546 510854
rect 329782 510618 329866 510854
rect 330102 510618 365546 510854
rect 365782 510618 365866 510854
rect 366102 510618 401546 510854
rect 401782 510618 401866 510854
rect 402102 510618 437546 510854
rect 437782 510618 437866 510854
rect 438102 510618 473546 510854
rect 473782 510618 473866 510854
rect 474102 510618 509546 510854
rect 509782 510618 509866 510854
rect 510102 510618 545546 510854
rect 545782 510618 545866 510854
rect 546102 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 587262 510854
rect 587498 510618 587582 510854
rect 587818 510618 588810 510854
rect -4886 510586 588810 510618
rect -2966 507454 586890 507486
rect -2966 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 109826 507454
rect 110062 507218 110146 507454
rect 110382 507218 145826 507454
rect 146062 507218 146146 507454
rect 146382 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 586890 507454
rect -2966 507134 586890 507218
rect -2966 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 109826 507134
rect 110062 506898 110146 507134
rect 110382 506898 145826 507134
rect 146062 506898 146146 507134
rect 146382 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 586890 507134
rect -2966 506866 586890 506898
rect -8726 500614 592650 500646
rect -8726 500378 -8694 500614
rect -8458 500378 -8374 500614
rect -8138 500378 30986 500614
rect 31222 500378 31306 500614
rect 31542 500378 66986 500614
rect 67222 500378 67306 500614
rect 67542 500378 102986 500614
rect 103222 500378 103306 500614
rect 103542 500378 138986 500614
rect 139222 500378 139306 500614
rect 139542 500378 426986 500614
rect 427222 500378 427306 500614
rect 427542 500378 462986 500614
rect 463222 500378 463306 500614
rect 463542 500378 498986 500614
rect 499222 500378 499306 500614
rect 499542 500378 534986 500614
rect 535222 500378 535306 500614
rect 535542 500378 570986 500614
rect 571222 500378 571306 500614
rect 571542 500378 592062 500614
rect 592298 500378 592382 500614
rect 592618 500378 592650 500614
rect -8726 500294 592650 500378
rect -8726 500058 -8694 500294
rect -8458 500058 -8374 500294
rect -8138 500058 30986 500294
rect 31222 500058 31306 500294
rect 31542 500058 66986 500294
rect 67222 500058 67306 500294
rect 67542 500058 102986 500294
rect 103222 500058 103306 500294
rect 103542 500058 138986 500294
rect 139222 500058 139306 500294
rect 139542 500058 426986 500294
rect 427222 500058 427306 500294
rect 427542 500058 462986 500294
rect 463222 500058 463306 500294
rect 463542 500058 498986 500294
rect 499222 500058 499306 500294
rect 499542 500058 534986 500294
rect 535222 500058 535306 500294
rect 535542 500058 570986 500294
rect 571222 500058 571306 500294
rect 571542 500058 592062 500294
rect 592298 500058 592382 500294
rect 592618 500058 592650 500294
rect -8726 500026 592650 500058
rect -6806 496894 590730 496926
rect -6806 496658 -6774 496894
rect -6538 496658 -6454 496894
rect -6218 496658 27266 496894
rect 27502 496658 27586 496894
rect 27822 496658 63266 496894
rect 63502 496658 63586 496894
rect 63822 496658 99266 496894
rect 99502 496658 99586 496894
rect 99822 496658 135266 496894
rect 135502 496658 135586 496894
rect 135822 496658 423266 496894
rect 423502 496658 423586 496894
rect 423822 496658 459266 496894
rect 459502 496658 459586 496894
rect 459822 496658 495266 496894
rect 495502 496658 495586 496894
rect 495822 496658 531266 496894
rect 531502 496658 531586 496894
rect 531822 496658 567266 496894
rect 567502 496658 567586 496894
rect 567822 496658 590142 496894
rect 590378 496658 590462 496894
rect 590698 496658 590730 496894
rect -6806 496574 590730 496658
rect -6806 496338 -6774 496574
rect -6538 496338 -6454 496574
rect -6218 496338 27266 496574
rect 27502 496338 27586 496574
rect 27822 496338 63266 496574
rect 63502 496338 63586 496574
rect 63822 496338 99266 496574
rect 99502 496338 99586 496574
rect 99822 496338 135266 496574
rect 135502 496338 135586 496574
rect 135822 496338 423266 496574
rect 423502 496338 423586 496574
rect 423822 496338 459266 496574
rect 459502 496338 459586 496574
rect 459822 496338 495266 496574
rect 495502 496338 495586 496574
rect 495822 496338 531266 496574
rect 531502 496338 531586 496574
rect 531822 496338 567266 496574
rect 567502 496338 567586 496574
rect 567822 496338 590142 496574
rect 590378 496338 590462 496574
rect 590698 496338 590730 496574
rect -6806 496306 590730 496338
rect -4886 493174 588810 493206
rect -4886 492938 -4854 493174
rect -4618 492938 -4534 493174
rect -4298 492938 23546 493174
rect 23782 492938 23866 493174
rect 24102 492938 59546 493174
rect 59782 492938 59866 493174
rect 60102 492938 95546 493174
rect 95782 492938 95866 493174
rect 96102 492938 131546 493174
rect 131782 492938 131866 493174
rect 132102 492938 455546 493174
rect 455782 492938 455866 493174
rect 456102 492938 491546 493174
rect 491782 492938 491866 493174
rect 492102 492938 527546 493174
rect 527782 492938 527866 493174
rect 528102 492938 563546 493174
rect 563782 492938 563866 493174
rect 564102 492938 588222 493174
rect 588458 492938 588542 493174
rect 588778 492938 588810 493174
rect -4886 492854 588810 492938
rect -4886 492618 -4854 492854
rect -4618 492618 -4534 492854
rect -4298 492618 23546 492854
rect 23782 492618 23866 492854
rect 24102 492618 59546 492854
rect 59782 492618 59866 492854
rect 60102 492618 95546 492854
rect 95782 492618 95866 492854
rect 96102 492618 131546 492854
rect 131782 492618 131866 492854
rect 132102 492618 455546 492854
rect 455782 492618 455866 492854
rect 456102 492618 491546 492854
rect 491782 492618 491866 492854
rect 492102 492618 527546 492854
rect 527782 492618 527866 492854
rect 528102 492618 563546 492854
rect 563782 492618 563866 492854
rect 564102 492618 588222 492854
rect 588458 492618 588542 492854
rect 588778 492618 588810 492854
rect -4886 492586 588810 492618
rect -2966 489454 586890 489486
rect -2966 489218 -2934 489454
rect -2698 489218 -2614 489454
rect -2378 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 91826 489454
rect 92062 489218 92146 489454
rect 92382 489218 127826 489454
rect 128062 489218 128146 489454
rect 128382 489218 185410 489454
rect 185646 489218 216130 489454
rect 216366 489218 246850 489454
rect 247086 489218 277570 489454
rect 277806 489218 308290 489454
rect 308526 489218 339010 489454
rect 339246 489218 369730 489454
rect 369966 489218 400450 489454
rect 400686 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 586302 489454
rect 586538 489218 586622 489454
rect 586858 489218 586890 489454
rect -2966 489134 586890 489218
rect -2966 488898 -2934 489134
rect -2698 488898 -2614 489134
rect -2378 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 91826 489134
rect 92062 488898 92146 489134
rect 92382 488898 127826 489134
rect 128062 488898 128146 489134
rect 128382 488898 185410 489134
rect 185646 488898 216130 489134
rect 216366 488898 246850 489134
rect 247086 488898 277570 489134
rect 277806 488898 308290 489134
rect 308526 488898 339010 489134
rect 339246 488898 369730 489134
rect 369966 488898 400450 489134
rect 400686 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 586302 489134
rect 586538 488898 586622 489134
rect 586858 488898 586890 489134
rect -2966 488866 586890 488898
rect -8726 482614 592650 482646
rect -8726 482378 -7734 482614
rect -7498 482378 -7414 482614
rect -7178 482378 12986 482614
rect 13222 482378 13306 482614
rect 13542 482378 48986 482614
rect 49222 482378 49306 482614
rect 49542 482378 84986 482614
rect 85222 482378 85306 482614
rect 85542 482378 120986 482614
rect 121222 482378 121306 482614
rect 121542 482378 156986 482614
rect 157222 482378 157306 482614
rect 157542 482378 444986 482614
rect 445222 482378 445306 482614
rect 445542 482378 480986 482614
rect 481222 482378 481306 482614
rect 481542 482378 516986 482614
rect 517222 482378 517306 482614
rect 517542 482378 552986 482614
rect 553222 482378 553306 482614
rect 553542 482378 591102 482614
rect 591338 482378 591422 482614
rect 591658 482378 592650 482614
rect -8726 482294 592650 482378
rect -8726 482058 -7734 482294
rect -7498 482058 -7414 482294
rect -7178 482058 12986 482294
rect 13222 482058 13306 482294
rect 13542 482058 48986 482294
rect 49222 482058 49306 482294
rect 49542 482058 84986 482294
rect 85222 482058 85306 482294
rect 85542 482058 120986 482294
rect 121222 482058 121306 482294
rect 121542 482058 156986 482294
rect 157222 482058 157306 482294
rect 157542 482058 444986 482294
rect 445222 482058 445306 482294
rect 445542 482058 480986 482294
rect 481222 482058 481306 482294
rect 481542 482058 516986 482294
rect 517222 482058 517306 482294
rect 517542 482058 552986 482294
rect 553222 482058 553306 482294
rect 553542 482058 591102 482294
rect 591338 482058 591422 482294
rect 591658 482058 592650 482294
rect -8726 482026 592650 482058
rect -6806 478894 590730 478926
rect -6806 478658 -5814 478894
rect -5578 478658 -5494 478894
rect -5258 478658 9266 478894
rect 9502 478658 9586 478894
rect 9822 478658 45266 478894
rect 45502 478658 45586 478894
rect 45822 478658 81266 478894
rect 81502 478658 81586 478894
rect 81822 478658 117266 478894
rect 117502 478658 117586 478894
rect 117822 478658 153266 478894
rect 153502 478658 153586 478894
rect 153822 478658 441266 478894
rect 441502 478658 441586 478894
rect 441822 478658 477266 478894
rect 477502 478658 477586 478894
rect 477822 478658 513266 478894
rect 513502 478658 513586 478894
rect 513822 478658 549266 478894
rect 549502 478658 549586 478894
rect 549822 478658 589182 478894
rect 589418 478658 589502 478894
rect 589738 478658 590730 478894
rect -6806 478574 590730 478658
rect -6806 478338 -5814 478574
rect -5578 478338 -5494 478574
rect -5258 478338 9266 478574
rect 9502 478338 9586 478574
rect 9822 478338 45266 478574
rect 45502 478338 45586 478574
rect 45822 478338 81266 478574
rect 81502 478338 81586 478574
rect 81822 478338 117266 478574
rect 117502 478338 117586 478574
rect 117822 478338 153266 478574
rect 153502 478338 153586 478574
rect 153822 478338 441266 478574
rect 441502 478338 441586 478574
rect 441822 478338 477266 478574
rect 477502 478338 477586 478574
rect 477822 478338 513266 478574
rect 513502 478338 513586 478574
rect 513822 478338 549266 478574
rect 549502 478338 549586 478574
rect 549822 478338 589182 478574
rect 589418 478338 589502 478574
rect 589738 478338 590730 478574
rect -6806 478306 590730 478338
rect -4886 475174 588810 475206
rect -4886 474938 -3894 475174
rect -3658 474938 -3574 475174
rect -3338 474938 5546 475174
rect 5782 474938 5866 475174
rect 6102 474938 41546 475174
rect 41782 474938 41866 475174
rect 42102 474938 77546 475174
rect 77782 474938 77866 475174
rect 78102 474938 113546 475174
rect 113782 474938 113866 475174
rect 114102 474938 149546 475174
rect 149782 474938 149866 475174
rect 150102 474938 437546 475174
rect 437782 474938 437866 475174
rect 438102 474938 473546 475174
rect 473782 474938 473866 475174
rect 474102 474938 509546 475174
rect 509782 474938 509866 475174
rect 510102 474938 545546 475174
rect 545782 474938 545866 475174
rect 546102 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 587262 475174
rect 587498 474938 587582 475174
rect 587818 474938 588810 475174
rect -4886 474854 588810 474938
rect -4886 474618 -3894 474854
rect -3658 474618 -3574 474854
rect -3338 474618 5546 474854
rect 5782 474618 5866 474854
rect 6102 474618 41546 474854
rect 41782 474618 41866 474854
rect 42102 474618 77546 474854
rect 77782 474618 77866 474854
rect 78102 474618 113546 474854
rect 113782 474618 113866 474854
rect 114102 474618 149546 474854
rect 149782 474618 149866 474854
rect 150102 474618 437546 474854
rect 437782 474618 437866 474854
rect 438102 474618 473546 474854
rect 473782 474618 473866 474854
rect 474102 474618 509546 474854
rect 509782 474618 509866 474854
rect 510102 474618 545546 474854
rect 545782 474618 545866 474854
rect 546102 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 587262 474854
rect 587498 474618 587582 474854
rect 587818 474618 588810 474854
rect -4886 474586 588810 474618
rect -2966 471454 586890 471486
rect -2966 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 170050 471454
rect 170286 471218 200770 471454
rect 201006 471218 231490 471454
rect 231726 471218 262210 471454
rect 262446 471218 292930 471454
rect 293166 471218 323650 471454
rect 323886 471218 354370 471454
rect 354606 471218 385090 471454
rect 385326 471218 415810 471454
rect 416046 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 586890 471454
rect -2966 471134 586890 471218
rect -2966 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 170050 471134
rect 170286 470898 200770 471134
rect 201006 470898 231490 471134
rect 231726 470898 262210 471134
rect 262446 470898 292930 471134
rect 293166 470898 323650 471134
rect 323886 470898 354370 471134
rect 354606 470898 385090 471134
rect 385326 470898 415810 471134
rect 416046 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 586890 471134
rect -2966 470866 586890 470898
rect -8726 464614 592650 464646
rect -8726 464378 -8694 464614
rect -8458 464378 -8374 464614
rect -8138 464378 30986 464614
rect 31222 464378 31306 464614
rect 31542 464378 66986 464614
rect 67222 464378 67306 464614
rect 67542 464378 102986 464614
rect 103222 464378 103306 464614
rect 103542 464378 138986 464614
rect 139222 464378 139306 464614
rect 139542 464378 426986 464614
rect 427222 464378 427306 464614
rect 427542 464378 462986 464614
rect 463222 464378 463306 464614
rect 463542 464378 498986 464614
rect 499222 464378 499306 464614
rect 499542 464378 534986 464614
rect 535222 464378 535306 464614
rect 535542 464378 570986 464614
rect 571222 464378 571306 464614
rect 571542 464378 592062 464614
rect 592298 464378 592382 464614
rect 592618 464378 592650 464614
rect -8726 464294 592650 464378
rect -8726 464058 -8694 464294
rect -8458 464058 -8374 464294
rect -8138 464058 30986 464294
rect 31222 464058 31306 464294
rect 31542 464058 66986 464294
rect 67222 464058 67306 464294
rect 67542 464058 102986 464294
rect 103222 464058 103306 464294
rect 103542 464058 138986 464294
rect 139222 464058 139306 464294
rect 139542 464058 426986 464294
rect 427222 464058 427306 464294
rect 427542 464058 462986 464294
rect 463222 464058 463306 464294
rect 463542 464058 498986 464294
rect 499222 464058 499306 464294
rect 499542 464058 534986 464294
rect 535222 464058 535306 464294
rect 535542 464058 570986 464294
rect 571222 464058 571306 464294
rect 571542 464058 592062 464294
rect 592298 464058 592382 464294
rect 592618 464058 592650 464294
rect -8726 464026 592650 464058
rect -6806 460894 590730 460926
rect -6806 460658 -6774 460894
rect -6538 460658 -6454 460894
rect -6218 460658 27266 460894
rect 27502 460658 27586 460894
rect 27822 460658 63266 460894
rect 63502 460658 63586 460894
rect 63822 460658 99266 460894
rect 99502 460658 99586 460894
rect 99822 460658 135266 460894
rect 135502 460658 135586 460894
rect 135822 460658 423266 460894
rect 423502 460658 423586 460894
rect 423822 460658 459266 460894
rect 459502 460658 459586 460894
rect 459822 460658 495266 460894
rect 495502 460658 495586 460894
rect 495822 460658 531266 460894
rect 531502 460658 531586 460894
rect 531822 460658 567266 460894
rect 567502 460658 567586 460894
rect 567822 460658 590142 460894
rect 590378 460658 590462 460894
rect 590698 460658 590730 460894
rect -6806 460574 590730 460658
rect -6806 460338 -6774 460574
rect -6538 460338 -6454 460574
rect -6218 460338 27266 460574
rect 27502 460338 27586 460574
rect 27822 460338 63266 460574
rect 63502 460338 63586 460574
rect 63822 460338 99266 460574
rect 99502 460338 99586 460574
rect 99822 460338 135266 460574
rect 135502 460338 135586 460574
rect 135822 460338 423266 460574
rect 423502 460338 423586 460574
rect 423822 460338 459266 460574
rect 459502 460338 459586 460574
rect 459822 460338 495266 460574
rect 495502 460338 495586 460574
rect 495822 460338 531266 460574
rect 531502 460338 531586 460574
rect 531822 460338 567266 460574
rect 567502 460338 567586 460574
rect 567822 460338 590142 460574
rect 590378 460338 590462 460574
rect 590698 460338 590730 460574
rect -6806 460306 590730 460338
rect -4886 457174 588810 457206
rect -4886 456938 -4854 457174
rect -4618 456938 -4534 457174
rect -4298 456938 23546 457174
rect 23782 456938 23866 457174
rect 24102 456938 59546 457174
rect 59782 456938 59866 457174
rect 60102 456938 95546 457174
rect 95782 456938 95866 457174
rect 96102 456938 131546 457174
rect 131782 456938 131866 457174
rect 132102 456938 455546 457174
rect 455782 456938 455866 457174
rect 456102 456938 491546 457174
rect 491782 456938 491866 457174
rect 492102 456938 527546 457174
rect 527782 456938 527866 457174
rect 528102 456938 563546 457174
rect 563782 456938 563866 457174
rect 564102 456938 588222 457174
rect 588458 456938 588542 457174
rect 588778 456938 588810 457174
rect -4886 456854 588810 456938
rect -4886 456618 -4854 456854
rect -4618 456618 -4534 456854
rect -4298 456618 23546 456854
rect 23782 456618 23866 456854
rect 24102 456618 59546 456854
rect 59782 456618 59866 456854
rect 60102 456618 95546 456854
rect 95782 456618 95866 456854
rect 96102 456618 131546 456854
rect 131782 456618 131866 456854
rect 132102 456618 455546 456854
rect 455782 456618 455866 456854
rect 456102 456618 491546 456854
rect 491782 456618 491866 456854
rect 492102 456618 527546 456854
rect 527782 456618 527866 456854
rect 528102 456618 563546 456854
rect 563782 456618 563866 456854
rect 564102 456618 588222 456854
rect 588458 456618 588542 456854
rect 588778 456618 588810 456854
rect -4886 456586 588810 456618
rect -2966 453454 586890 453486
rect -2966 453218 -2934 453454
rect -2698 453218 -2614 453454
rect -2378 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 91826 453454
rect 92062 453218 92146 453454
rect 92382 453218 127826 453454
rect 128062 453218 128146 453454
rect 128382 453218 185410 453454
rect 185646 453218 216130 453454
rect 216366 453218 246850 453454
rect 247086 453218 277570 453454
rect 277806 453218 308290 453454
rect 308526 453218 339010 453454
rect 339246 453218 369730 453454
rect 369966 453218 400450 453454
rect 400686 453218 451826 453454
rect 452062 453218 452146 453454
rect 452382 453218 487826 453454
rect 488062 453218 488146 453454
rect 488382 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 586302 453454
rect 586538 453218 586622 453454
rect 586858 453218 586890 453454
rect -2966 453134 586890 453218
rect -2966 452898 -2934 453134
rect -2698 452898 -2614 453134
rect -2378 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 91826 453134
rect 92062 452898 92146 453134
rect 92382 452898 127826 453134
rect 128062 452898 128146 453134
rect 128382 452898 185410 453134
rect 185646 452898 216130 453134
rect 216366 452898 246850 453134
rect 247086 452898 277570 453134
rect 277806 452898 308290 453134
rect 308526 452898 339010 453134
rect 339246 452898 369730 453134
rect 369966 452898 400450 453134
rect 400686 452898 451826 453134
rect 452062 452898 452146 453134
rect 452382 452898 487826 453134
rect 488062 452898 488146 453134
rect 488382 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 586302 453134
rect 586538 452898 586622 453134
rect 586858 452898 586890 453134
rect -2966 452866 586890 452898
rect -8726 446614 592650 446646
rect -8726 446378 -7734 446614
rect -7498 446378 -7414 446614
rect -7178 446378 12986 446614
rect 13222 446378 13306 446614
rect 13542 446378 48986 446614
rect 49222 446378 49306 446614
rect 49542 446378 84986 446614
rect 85222 446378 85306 446614
rect 85542 446378 120986 446614
rect 121222 446378 121306 446614
rect 121542 446378 156986 446614
rect 157222 446378 157306 446614
rect 157542 446378 444986 446614
rect 445222 446378 445306 446614
rect 445542 446378 480986 446614
rect 481222 446378 481306 446614
rect 481542 446378 516986 446614
rect 517222 446378 517306 446614
rect 517542 446378 552986 446614
rect 553222 446378 553306 446614
rect 553542 446378 591102 446614
rect 591338 446378 591422 446614
rect 591658 446378 592650 446614
rect -8726 446294 592650 446378
rect -8726 446058 -7734 446294
rect -7498 446058 -7414 446294
rect -7178 446058 12986 446294
rect 13222 446058 13306 446294
rect 13542 446058 48986 446294
rect 49222 446058 49306 446294
rect 49542 446058 84986 446294
rect 85222 446058 85306 446294
rect 85542 446058 120986 446294
rect 121222 446058 121306 446294
rect 121542 446058 156986 446294
rect 157222 446058 157306 446294
rect 157542 446058 444986 446294
rect 445222 446058 445306 446294
rect 445542 446058 480986 446294
rect 481222 446058 481306 446294
rect 481542 446058 516986 446294
rect 517222 446058 517306 446294
rect 517542 446058 552986 446294
rect 553222 446058 553306 446294
rect 553542 446058 591102 446294
rect 591338 446058 591422 446294
rect 591658 446058 592650 446294
rect -8726 446026 592650 446058
rect -6806 442894 590730 442926
rect -6806 442658 -5814 442894
rect -5578 442658 -5494 442894
rect -5258 442658 9266 442894
rect 9502 442658 9586 442894
rect 9822 442658 45266 442894
rect 45502 442658 45586 442894
rect 45822 442658 81266 442894
rect 81502 442658 81586 442894
rect 81822 442658 117266 442894
rect 117502 442658 117586 442894
rect 117822 442658 153266 442894
rect 153502 442658 153586 442894
rect 153822 442658 441266 442894
rect 441502 442658 441586 442894
rect 441822 442658 477266 442894
rect 477502 442658 477586 442894
rect 477822 442658 513266 442894
rect 513502 442658 513586 442894
rect 513822 442658 549266 442894
rect 549502 442658 549586 442894
rect 549822 442658 589182 442894
rect 589418 442658 589502 442894
rect 589738 442658 590730 442894
rect -6806 442574 590730 442658
rect -6806 442338 -5814 442574
rect -5578 442338 -5494 442574
rect -5258 442338 9266 442574
rect 9502 442338 9586 442574
rect 9822 442338 45266 442574
rect 45502 442338 45586 442574
rect 45822 442338 81266 442574
rect 81502 442338 81586 442574
rect 81822 442338 117266 442574
rect 117502 442338 117586 442574
rect 117822 442338 153266 442574
rect 153502 442338 153586 442574
rect 153822 442338 441266 442574
rect 441502 442338 441586 442574
rect 441822 442338 477266 442574
rect 477502 442338 477586 442574
rect 477822 442338 513266 442574
rect 513502 442338 513586 442574
rect 513822 442338 549266 442574
rect 549502 442338 549586 442574
rect 549822 442338 589182 442574
rect 589418 442338 589502 442574
rect 589738 442338 590730 442574
rect -6806 442306 590730 442338
rect -4886 439174 588810 439206
rect -4886 438938 -3894 439174
rect -3658 438938 -3574 439174
rect -3338 438938 5546 439174
rect 5782 438938 5866 439174
rect 6102 438938 41546 439174
rect 41782 438938 41866 439174
rect 42102 438938 77546 439174
rect 77782 438938 77866 439174
rect 78102 438938 113546 439174
rect 113782 438938 113866 439174
rect 114102 438938 149546 439174
rect 149782 438938 149866 439174
rect 150102 438938 437546 439174
rect 437782 438938 437866 439174
rect 438102 438938 473546 439174
rect 473782 438938 473866 439174
rect 474102 438938 509546 439174
rect 509782 438938 509866 439174
rect 510102 438938 545546 439174
rect 545782 438938 545866 439174
rect 546102 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 587262 439174
rect 587498 438938 587582 439174
rect 587818 438938 588810 439174
rect -4886 438854 588810 438938
rect -4886 438618 -3894 438854
rect -3658 438618 -3574 438854
rect -3338 438618 5546 438854
rect 5782 438618 5866 438854
rect 6102 438618 41546 438854
rect 41782 438618 41866 438854
rect 42102 438618 77546 438854
rect 77782 438618 77866 438854
rect 78102 438618 113546 438854
rect 113782 438618 113866 438854
rect 114102 438618 149546 438854
rect 149782 438618 149866 438854
rect 150102 438618 437546 438854
rect 437782 438618 437866 438854
rect 438102 438618 473546 438854
rect 473782 438618 473866 438854
rect 474102 438618 509546 438854
rect 509782 438618 509866 438854
rect 510102 438618 545546 438854
rect 545782 438618 545866 438854
rect 546102 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 587262 438854
rect 587498 438618 587582 438854
rect 587818 438618 588810 438854
rect -4886 438586 588810 438618
rect -2966 435454 586890 435486
rect -2966 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 73826 435454
rect 74062 435218 74146 435454
rect 74382 435218 109826 435454
rect 110062 435218 110146 435454
rect 110382 435218 145826 435454
rect 146062 435218 146146 435454
rect 146382 435218 170050 435454
rect 170286 435218 200770 435454
rect 201006 435218 231490 435454
rect 231726 435218 262210 435454
rect 262446 435218 292930 435454
rect 293166 435218 323650 435454
rect 323886 435218 354370 435454
rect 354606 435218 385090 435454
rect 385326 435218 415810 435454
rect 416046 435218 433826 435454
rect 434062 435218 434146 435454
rect 434382 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 586890 435454
rect -2966 435134 586890 435218
rect -2966 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 73826 435134
rect 74062 434898 74146 435134
rect 74382 434898 109826 435134
rect 110062 434898 110146 435134
rect 110382 434898 145826 435134
rect 146062 434898 146146 435134
rect 146382 434898 170050 435134
rect 170286 434898 200770 435134
rect 201006 434898 231490 435134
rect 231726 434898 262210 435134
rect 262446 434898 292930 435134
rect 293166 434898 323650 435134
rect 323886 434898 354370 435134
rect 354606 434898 385090 435134
rect 385326 434898 415810 435134
rect 416046 434898 433826 435134
rect 434062 434898 434146 435134
rect 434382 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 586890 435134
rect -2966 434866 586890 434898
rect -8726 428614 592650 428646
rect -8726 428378 -8694 428614
rect -8458 428378 -8374 428614
rect -8138 428378 30986 428614
rect 31222 428378 31306 428614
rect 31542 428378 66986 428614
rect 67222 428378 67306 428614
rect 67542 428378 102986 428614
rect 103222 428378 103306 428614
rect 103542 428378 138986 428614
rect 139222 428378 139306 428614
rect 139542 428378 426986 428614
rect 427222 428378 427306 428614
rect 427542 428378 462986 428614
rect 463222 428378 463306 428614
rect 463542 428378 498986 428614
rect 499222 428378 499306 428614
rect 499542 428378 534986 428614
rect 535222 428378 535306 428614
rect 535542 428378 570986 428614
rect 571222 428378 571306 428614
rect 571542 428378 592062 428614
rect 592298 428378 592382 428614
rect 592618 428378 592650 428614
rect -8726 428294 592650 428378
rect -8726 428058 -8694 428294
rect -8458 428058 -8374 428294
rect -8138 428058 30986 428294
rect 31222 428058 31306 428294
rect 31542 428058 66986 428294
rect 67222 428058 67306 428294
rect 67542 428058 102986 428294
rect 103222 428058 103306 428294
rect 103542 428058 138986 428294
rect 139222 428058 139306 428294
rect 139542 428058 426986 428294
rect 427222 428058 427306 428294
rect 427542 428058 462986 428294
rect 463222 428058 463306 428294
rect 463542 428058 498986 428294
rect 499222 428058 499306 428294
rect 499542 428058 534986 428294
rect 535222 428058 535306 428294
rect 535542 428058 570986 428294
rect 571222 428058 571306 428294
rect 571542 428058 592062 428294
rect 592298 428058 592382 428294
rect 592618 428058 592650 428294
rect -8726 428026 592650 428058
rect -6806 424894 590730 424926
rect -6806 424658 -6774 424894
rect -6538 424658 -6454 424894
rect -6218 424658 27266 424894
rect 27502 424658 27586 424894
rect 27822 424658 63266 424894
rect 63502 424658 63586 424894
rect 63822 424658 99266 424894
rect 99502 424658 99586 424894
rect 99822 424658 135266 424894
rect 135502 424658 135586 424894
rect 135822 424658 423266 424894
rect 423502 424658 423586 424894
rect 423822 424658 459266 424894
rect 459502 424658 459586 424894
rect 459822 424658 495266 424894
rect 495502 424658 495586 424894
rect 495822 424658 531266 424894
rect 531502 424658 531586 424894
rect 531822 424658 567266 424894
rect 567502 424658 567586 424894
rect 567822 424658 590142 424894
rect 590378 424658 590462 424894
rect 590698 424658 590730 424894
rect -6806 424574 590730 424658
rect -6806 424338 -6774 424574
rect -6538 424338 -6454 424574
rect -6218 424338 27266 424574
rect 27502 424338 27586 424574
rect 27822 424338 63266 424574
rect 63502 424338 63586 424574
rect 63822 424338 99266 424574
rect 99502 424338 99586 424574
rect 99822 424338 135266 424574
rect 135502 424338 135586 424574
rect 135822 424338 423266 424574
rect 423502 424338 423586 424574
rect 423822 424338 459266 424574
rect 459502 424338 459586 424574
rect 459822 424338 495266 424574
rect 495502 424338 495586 424574
rect 495822 424338 531266 424574
rect 531502 424338 531586 424574
rect 531822 424338 567266 424574
rect 567502 424338 567586 424574
rect 567822 424338 590142 424574
rect 590378 424338 590462 424574
rect 590698 424338 590730 424574
rect -6806 424306 590730 424338
rect -4886 421174 588810 421206
rect -4886 420938 -4854 421174
rect -4618 420938 -4534 421174
rect -4298 420938 23546 421174
rect 23782 420938 23866 421174
rect 24102 420938 59546 421174
rect 59782 420938 59866 421174
rect 60102 420938 95546 421174
rect 95782 420938 95866 421174
rect 96102 420938 131546 421174
rect 131782 420938 131866 421174
rect 132102 420938 455546 421174
rect 455782 420938 455866 421174
rect 456102 420938 491546 421174
rect 491782 420938 491866 421174
rect 492102 420938 527546 421174
rect 527782 420938 527866 421174
rect 528102 420938 563546 421174
rect 563782 420938 563866 421174
rect 564102 420938 588222 421174
rect 588458 420938 588542 421174
rect 588778 420938 588810 421174
rect -4886 420854 588810 420938
rect -4886 420618 -4854 420854
rect -4618 420618 -4534 420854
rect -4298 420618 23546 420854
rect 23782 420618 23866 420854
rect 24102 420618 59546 420854
rect 59782 420618 59866 420854
rect 60102 420618 95546 420854
rect 95782 420618 95866 420854
rect 96102 420618 131546 420854
rect 131782 420618 131866 420854
rect 132102 420618 455546 420854
rect 455782 420618 455866 420854
rect 456102 420618 491546 420854
rect 491782 420618 491866 420854
rect 492102 420618 527546 420854
rect 527782 420618 527866 420854
rect 528102 420618 563546 420854
rect 563782 420618 563866 420854
rect 564102 420618 588222 420854
rect 588458 420618 588542 420854
rect 588778 420618 588810 420854
rect -4886 420586 588810 420618
rect -2966 417454 586890 417486
rect -2966 417218 -2934 417454
rect -2698 417218 -2614 417454
rect -2378 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 91826 417454
rect 92062 417218 92146 417454
rect 92382 417218 127826 417454
rect 128062 417218 128146 417454
rect 128382 417218 185410 417454
rect 185646 417218 216130 417454
rect 216366 417218 246850 417454
rect 247086 417218 277570 417454
rect 277806 417218 308290 417454
rect 308526 417218 339010 417454
rect 339246 417218 369730 417454
rect 369966 417218 400450 417454
rect 400686 417218 451826 417454
rect 452062 417218 452146 417454
rect 452382 417218 487826 417454
rect 488062 417218 488146 417454
rect 488382 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 586302 417454
rect 586538 417218 586622 417454
rect 586858 417218 586890 417454
rect -2966 417134 586890 417218
rect -2966 416898 -2934 417134
rect -2698 416898 -2614 417134
rect -2378 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 91826 417134
rect 92062 416898 92146 417134
rect 92382 416898 127826 417134
rect 128062 416898 128146 417134
rect 128382 416898 185410 417134
rect 185646 416898 216130 417134
rect 216366 416898 246850 417134
rect 247086 416898 277570 417134
rect 277806 416898 308290 417134
rect 308526 416898 339010 417134
rect 339246 416898 369730 417134
rect 369966 416898 400450 417134
rect 400686 416898 451826 417134
rect 452062 416898 452146 417134
rect 452382 416898 487826 417134
rect 488062 416898 488146 417134
rect 488382 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 586302 417134
rect 586538 416898 586622 417134
rect 586858 416898 586890 417134
rect -2966 416866 586890 416898
rect -8726 410614 592650 410646
rect -8726 410378 -7734 410614
rect -7498 410378 -7414 410614
rect -7178 410378 12986 410614
rect 13222 410378 13306 410614
rect 13542 410378 48986 410614
rect 49222 410378 49306 410614
rect 49542 410378 84986 410614
rect 85222 410378 85306 410614
rect 85542 410378 120986 410614
rect 121222 410378 121306 410614
rect 121542 410378 156986 410614
rect 157222 410378 157306 410614
rect 157542 410378 444986 410614
rect 445222 410378 445306 410614
rect 445542 410378 480986 410614
rect 481222 410378 481306 410614
rect 481542 410378 516986 410614
rect 517222 410378 517306 410614
rect 517542 410378 552986 410614
rect 553222 410378 553306 410614
rect 553542 410378 591102 410614
rect 591338 410378 591422 410614
rect 591658 410378 592650 410614
rect -8726 410294 592650 410378
rect -8726 410058 -7734 410294
rect -7498 410058 -7414 410294
rect -7178 410058 12986 410294
rect 13222 410058 13306 410294
rect 13542 410058 48986 410294
rect 49222 410058 49306 410294
rect 49542 410058 84986 410294
rect 85222 410058 85306 410294
rect 85542 410058 120986 410294
rect 121222 410058 121306 410294
rect 121542 410058 156986 410294
rect 157222 410058 157306 410294
rect 157542 410058 444986 410294
rect 445222 410058 445306 410294
rect 445542 410058 480986 410294
rect 481222 410058 481306 410294
rect 481542 410058 516986 410294
rect 517222 410058 517306 410294
rect 517542 410058 552986 410294
rect 553222 410058 553306 410294
rect 553542 410058 591102 410294
rect 591338 410058 591422 410294
rect 591658 410058 592650 410294
rect -8726 410026 592650 410058
rect -6806 406894 590730 406926
rect -6806 406658 -5814 406894
rect -5578 406658 -5494 406894
rect -5258 406658 9266 406894
rect 9502 406658 9586 406894
rect 9822 406658 45266 406894
rect 45502 406658 45586 406894
rect 45822 406658 81266 406894
rect 81502 406658 81586 406894
rect 81822 406658 117266 406894
rect 117502 406658 117586 406894
rect 117822 406658 153266 406894
rect 153502 406658 153586 406894
rect 153822 406658 441266 406894
rect 441502 406658 441586 406894
rect 441822 406658 477266 406894
rect 477502 406658 477586 406894
rect 477822 406658 513266 406894
rect 513502 406658 513586 406894
rect 513822 406658 549266 406894
rect 549502 406658 549586 406894
rect 549822 406658 589182 406894
rect 589418 406658 589502 406894
rect 589738 406658 590730 406894
rect -6806 406574 590730 406658
rect -6806 406338 -5814 406574
rect -5578 406338 -5494 406574
rect -5258 406338 9266 406574
rect 9502 406338 9586 406574
rect 9822 406338 45266 406574
rect 45502 406338 45586 406574
rect 45822 406338 81266 406574
rect 81502 406338 81586 406574
rect 81822 406338 117266 406574
rect 117502 406338 117586 406574
rect 117822 406338 153266 406574
rect 153502 406338 153586 406574
rect 153822 406338 441266 406574
rect 441502 406338 441586 406574
rect 441822 406338 477266 406574
rect 477502 406338 477586 406574
rect 477822 406338 513266 406574
rect 513502 406338 513586 406574
rect 513822 406338 549266 406574
rect 549502 406338 549586 406574
rect 549822 406338 589182 406574
rect 589418 406338 589502 406574
rect 589738 406338 590730 406574
rect -6806 406306 590730 406338
rect -4886 403174 588810 403206
rect -4886 402938 -3894 403174
rect -3658 402938 -3574 403174
rect -3338 402938 5546 403174
rect 5782 402938 5866 403174
rect 6102 402938 41546 403174
rect 41782 402938 41866 403174
rect 42102 402938 77546 403174
rect 77782 402938 77866 403174
rect 78102 402938 113546 403174
rect 113782 402938 113866 403174
rect 114102 402938 149546 403174
rect 149782 402938 149866 403174
rect 150102 402938 437546 403174
rect 437782 402938 437866 403174
rect 438102 402938 473546 403174
rect 473782 402938 473866 403174
rect 474102 402938 509546 403174
rect 509782 402938 509866 403174
rect 510102 402938 545546 403174
rect 545782 402938 545866 403174
rect 546102 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 587262 403174
rect 587498 402938 587582 403174
rect 587818 402938 588810 403174
rect -4886 402854 588810 402938
rect -4886 402618 -3894 402854
rect -3658 402618 -3574 402854
rect -3338 402618 5546 402854
rect 5782 402618 5866 402854
rect 6102 402618 41546 402854
rect 41782 402618 41866 402854
rect 42102 402618 77546 402854
rect 77782 402618 77866 402854
rect 78102 402618 113546 402854
rect 113782 402618 113866 402854
rect 114102 402618 149546 402854
rect 149782 402618 149866 402854
rect 150102 402618 437546 402854
rect 437782 402618 437866 402854
rect 438102 402618 473546 402854
rect 473782 402618 473866 402854
rect 474102 402618 509546 402854
rect 509782 402618 509866 402854
rect 510102 402618 545546 402854
rect 545782 402618 545866 402854
rect 546102 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 587262 402854
rect 587498 402618 587582 402854
rect 587818 402618 588810 402854
rect -4886 402586 588810 402618
rect -2966 399454 586890 399486
rect -2966 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 73826 399454
rect 74062 399218 74146 399454
rect 74382 399218 109826 399454
rect 110062 399218 110146 399454
rect 110382 399218 145826 399454
rect 146062 399218 146146 399454
rect 146382 399218 170050 399454
rect 170286 399218 200770 399454
rect 201006 399218 231490 399454
rect 231726 399218 262210 399454
rect 262446 399218 292930 399454
rect 293166 399218 323650 399454
rect 323886 399218 354370 399454
rect 354606 399218 385090 399454
rect 385326 399218 415810 399454
rect 416046 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 586890 399454
rect -2966 399134 586890 399218
rect -2966 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 73826 399134
rect 74062 398898 74146 399134
rect 74382 398898 109826 399134
rect 110062 398898 110146 399134
rect 110382 398898 145826 399134
rect 146062 398898 146146 399134
rect 146382 398898 170050 399134
rect 170286 398898 200770 399134
rect 201006 398898 231490 399134
rect 231726 398898 262210 399134
rect 262446 398898 292930 399134
rect 293166 398898 323650 399134
rect 323886 398898 354370 399134
rect 354606 398898 385090 399134
rect 385326 398898 415810 399134
rect 416046 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 586890 399134
rect -2966 398866 586890 398898
rect -8726 392614 592650 392646
rect -8726 392378 -8694 392614
rect -8458 392378 -8374 392614
rect -8138 392378 30986 392614
rect 31222 392378 31306 392614
rect 31542 392378 66986 392614
rect 67222 392378 67306 392614
rect 67542 392378 102986 392614
rect 103222 392378 103306 392614
rect 103542 392378 138986 392614
rect 139222 392378 139306 392614
rect 139542 392378 426986 392614
rect 427222 392378 427306 392614
rect 427542 392378 462986 392614
rect 463222 392378 463306 392614
rect 463542 392378 498986 392614
rect 499222 392378 499306 392614
rect 499542 392378 534986 392614
rect 535222 392378 535306 392614
rect 535542 392378 570986 392614
rect 571222 392378 571306 392614
rect 571542 392378 592062 392614
rect 592298 392378 592382 392614
rect 592618 392378 592650 392614
rect -8726 392294 592650 392378
rect -8726 392058 -8694 392294
rect -8458 392058 -8374 392294
rect -8138 392058 30986 392294
rect 31222 392058 31306 392294
rect 31542 392058 66986 392294
rect 67222 392058 67306 392294
rect 67542 392058 102986 392294
rect 103222 392058 103306 392294
rect 103542 392058 138986 392294
rect 139222 392058 139306 392294
rect 139542 392058 426986 392294
rect 427222 392058 427306 392294
rect 427542 392058 462986 392294
rect 463222 392058 463306 392294
rect 463542 392058 498986 392294
rect 499222 392058 499306 392294
rect 499542 392058 534986 392294
rect 535222 392058 535306 392294
rect 535542 392058 570986 392294
rect 571222 392058 571306 392294
rect 571542 392058 592062 392294
rect 592298 392058 592382 392294
rect 592618 392058 592650 392294
rect -8726 392026 592650 392058
rect -6806 388894 590730 388926
rect -6806 388658 -6774 388894
rect -6538 388658 -6454 388894
rect -6218 388658 27266 388894
rect 27502 388658 27586 388894
rect 27822 388658 63266 388894
rect 63502 388658 63586 388894
rect 63822 388658 99266 388894
rect 99502 388658 99586 388894
rect 99822 388658 135266 388894
rect 135502 388658 135586 388894
rect 135822 388658 423266 388894
rect 423502 388658 423586 388894
rect 423822 388658 459266 388894
rect 459502 388658 459586 388894
rect 459822 388658 495266 388894
rect 495502 388658 495586 388894
rect 495822 388658 531266 388894
rect 531502 388658 531586 388894
rect 531822 388658 567266 388894
rect 567502 388658 567586 388894
rect 567822 388658 590142 388894
rect 590378 388658 590462 388894
rect 590698 388658 590730 388894
rect -6806 388574 590730 388658
rect -6806 388338 -6774 388574
rect -6538 388338 -6454 388574
rect -6218 388338 27266 388574
rect 27502 388338 27586 388574
rect 27822 388338 63266 388574
rect 63502 388338 63586 388574
rect 63822 388338 99266 388574
rect 99502 388338 99586 388574
rect 99822 388338 135266 388574
rect 135502 388338 135586 388574
rect 135822 388338 423266 388574
rect 423502 388338 423586 388574
rect 423822 388338 459266 388574
rect 459502 388338 459586 388574
rect 459822 388338 495266 388574
rect 495502 388338 495586 388574
rect 495822 388338 531266 388574
rect 531502 388338 531586 388574
rect 531822 388338 567266 388574
rect 567502 388338 567586 388574
rect 567822 388338 590142 388574
rect 590378 388338 590462 388574
rect 590698 388338 590730 388574
rect -6806 388306 590730 388338
rect -4886 385174 588810 385206
rect -4886 384938 -4854 385174
rect -4618 384938 -4534 385174
rect -4298 384938 23546 385174
rect 23782 384938 23866 385174
rect 24102 384938 59546 385174
rect 59782 384938 59866 385174
rect 60102 384938 95546 385174
rect 95782 384938 95866 385174
rect 96102 384938 131546 385174
rect 131782 384938 131866 385174
rect 132102 384938 455546 385174
rect 455782 384938 455866 385174
rect 456102 384938 491546 385174
rect 491782 384938 491866 385174
rect 492102 384938 527546 385174
rect 527782 384938 527866 385174
rect 528102 384938 563546 385174
rect 563782 384938 563866 385174
rect 564102 384938 588222 385174
rect 588458 384938 588542 385174
rect 588778 384938 588810 385174
rect -4886 384854 588810 384938
rect -4886 384618 -4854 384854
rect -4618 384618 -4534 384854
rect -4298 384618 23546 384854
rect 23782 384618 23866 384854
rect 24102 384618 59546 384854
rect 59782 384618 59866 384854
rect 60102 384618 95546 384854
rect 95782 384618 95866 384854
rect 96102 384618 131546 384854
rect 131782 384618 131866 384854
rect 132102 384618 455546 384854
rect 455782 384618 455866 384854
rect 456102 384618 491546 384854
rect 491782 384618 491866 384854
rect 492102 384618 527546 384854
rect 527782 384618 527866 384854
rect 528102 384618 563546 384854
rect 563782 384618 563866 384854
rect 564102 384618 588222 384854
rect 588458 384618 588542 384854
rect 588778 384618 588810 384854
rect -4886 384586 588810 384618
rect -2966 381454 586890 381486
rect -2966 381218 -2934 381454
rect -2698 381218 -2614 381454
rect -2378 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 91826 381454
rect 92062 381218 92146 381454
rect 92382 381218 127826 381454
rect 128062 381218 128146 381454
rect 128382 381218 185410 381454
rect 185646 381218 216130 381454
rect 216366 381218 246850 381454
rect 247086 381218 277570 381454
rect 277806 381218 308290 381454
rect 308526 381218 339010 381454
rect 339246 381218 369730 381454
rect 369966 381218 400450 381454
rect 400686 381218 451826 381454
rect 452062 381218 452146 381454
rect 452382 381218 487826 381454
rect 488062 381218 488146 381454
rect 488382 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 586302 381454
rect 586538 381218 586622 381454
rect 586858 381218 586890 381454
rect -2966 381134 586890 381218
rect -2966 380898 -2934 381134
rect -2698 380898 -2614 381134
rect -2378 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 91826 381134
rect 92062 380898 92146 381134
rect 92382 380898 127826 381134
rect 128062 380898 128146 381134
rect 128382 380898 185410 381134
rect 185646 380898 216130 381134
rect 216366 380898 246850 381134
rect 247086 380898 277570 381134
rect 277806 380898 308290 381134
rect 308526 380898 339010 381134
rect 339246 380898 369730 381134
rect 369966 380898 400450 381134
rect 400686 380898 451826 381134
rect 452062 380898 452146 381134
rect 452382 380898 487826 381134
rect 488062 380898 488146 381134
rect 488382 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 586302 381134
rect 586538 380898 586622 381134
rect 586858 380898 586890 381134
rect -2966 380866 586890 380898
rect -8726 374614 592650 374646
rect -8726 374378 -7734 374614
rect -7498 374378 -7414 374614
rect -7178 374378 12986 374614
rect 13222 374378 13306 374614
rect 13542 374378 48986 374614
rect 49222 374378 49306 374614
rect 49542 374378 84986 374614
rect 85222 374378 85306 374614
rect 85542 374378 120986 374614
rect 121222 374378 121306 374614
rect 121542 374378 156986 374614
rect 157222 374378 157306 374614
rect 157542 374378 444986 374614
rect 445222 374378 445306 374614
rect 445542 374378 480986 374614
rect 481222 374378 481306 374614
rect 481542 374378 516986 374614
rect 517222 374378 517306 374614
rect 517542 374378 552986 374614
rect 553222 374378 553306 374614
rect 553542 374378 591102 374614
rect 591338 374378 591422 374614
rect 591658 374378 592650 374614
rect -8726 374294 592650 374378
rect -8726 374058 -7734 374294
rect -7498 374058 -7414 374294
rect -7178 374058 12986 374294
rect 13222 374058 13306 374294
rect 13542 374058 48986 374294
rect 49222 374058 49306 374294
rect 49542 374058 84986 374294
rect 85222 374058 85306 374294
rect 85542 374058 120986 374294
rect 121222 374058 121306 374294
rect 121542 374058 156986 374294
rect 157222 374058 157306 374294
rect 157542 374058 444986 374294
rect 445222 374058 445306 374294
rect 445542 374058 480986 374294
rect 481222 374058 481306 374294
rect 481542 374058 516986 374294
rect 517222 374058 517306 374294
rect 517542 374058 552986 374294
rect 553222 374058 553306 374294
rect 553542 374058 591102 374294
rect 591338 374058 591422 374294
rect 591658 374058 592650 374294
rect -8726 374026 592650 374058
rect -6806 370894 590730 370926
rect -6806 370658 -5814 370894
rect -5578 370658 -5494 370894
rect -5258 370658 9266 370894
rect 9502 370658 9586 370894
rect 9822 370658 45266 370894
rect 45502 370658 45586 370894
rect 45822 370658 81266 370894
rect 81502 370658 81586 370894
rect 81822 370658 117266 370894
rect 117502 370658 117586 370894
rect 117822 370658 153266 370894
rect 153502 370658 153586 370894
rect 153822 370658 441266 370894
rect 441502 370658 441586 370894
rect 441822 370658 477266 370894
rect 477502 370658 477586 370894
rect 477822 370658 513266 370894
rect 513502 370658 513586 370894
rect 513822 370658 549266 370894
rect 549502 370658 549586 370894
rect 549822 370658 589182 370894
rect 589418 370658 589502 370894
rect 589738 370658 590730 370894
rect -6806 370574 590730 370658
rect -6806 370338 -5814 370574
rect -5578 370338 -5494 370574
rect -5258 370338 9266 370574
rect 9502 370338 9586 370574
rect 9822 370338 45266 370574
rect 45502 370338 45586 370574
rect 45822 370338 81266 370574
rect 81502 370338 81586 370574
rect 81822 370338 117266 370574
rect 117502 370338 117586 370574
rect 117822 370338 153266 370574
rect 153502 370338 153586 370574
rect 153822 370338 441266 370574
rect 441502 370338 441586 370574
rect 441822 370338 477266 370574
rect 477502 370338 477586 370574
rect 477822 370338 513266 370574
rect 513502 370338 513586 370574
rect 513822 370338 549266 370574
rect 549502 370338 549586 370574
rect 549822 370338 589182 370574
rect 589418 370338 589502 370574
rect 589738 370338 590730 370574
rect -6806 370306 590730 370338
rect -4886 367174 588810 367206
rect -4886 366938 -3894 367174
rect -3658 366938 -3574 367174
rect -3338 366938 5546 367174
rect 5782 366938 5866 367174
rect 6102 366938 41546 367174
rect 41782 366938 41866 367174
rect 42102 366938 77546 367174
rect 77782 366938 77866 367174
rect 78102 366938 113546 367174
rect 113782 366938 113866 367174
rect 114102 366938 149546 367174
rect 149782 366938 149866 367174
rect 150102 366938 437546 367174
rect 437782 366938 437866 367174
rect 438102 366938 473546 367174
rect 473782 366938 473866 367174
rect 474102 366938 509546 367174
rect 509782 366938 509866 367174
rect 510102 366938 545546 367174
rect 545782 366938 545866 367174
rect 546102 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 587262 367174
rect 587498 366938 587582 367174
rect 587818 366938 588810 367174
rect -4886 366854 588810 366938
rect -4886 366618 -3894 366854
rect -3658 366618 -3574 366854
rect -3338 366618 5546 366854
rect 5782 366618 5866 366854
rect 6102 366618 41546 366854
rect 41782 366618 41866 366854
rect 42102 366618 77546 366854
rect 77782 366618 77866 366854
rect 78102 366618 113546 366854
rect 113782 366618 113866 366854
rect 114102 366618 149546 366854
rect 149782 366618 149866 366854
rect 150102 366618 437546 366854
rect 437782 366618 437866 366854
rect 438102 366618 473546 366854
rect 473782 366618 473866 366854
rect 474102 366618 509546 366854
rect 509782 366618 509866 366854
rect 510102 366618 545546 366854
rect 545782 366618 545866 366854
rect 546102 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 587262 366854
rect 587498 366618 587582 366854
rect 587818 366618 588810 366854
rect -4886 366586 588810 366618
rect -2966 363454 586890 363486
rect -2966 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 109826 363454
rect 110062 363218 110146 363454
rect 110382 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 170050 363454
rect 170286 363218 200770 363454
rect 201006 363218 231490 363454
rect 231726 363218 262210 363454
rect 262446 363218 292930 363454
rect 293166 363218 323650 363454
rect 323886 363218 354370 363454
rect 354606 363218 385090 363454
rect 385326 363218 415810 363454
rect 416046 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 586890 363454
rect -2966 363134 586890 363218
rect -2966 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 109826 363134
rect 110062 362898 110146 363134
rect 110382 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 170050 363134
rect 170286 362898 200770 363134
rect 201006 362898 231490 363134
rect 231726 362898 262210 363134
rect 262446 362898 292930 363134
rect 293166 362898 323650 363134
rect 323886 362898 354370 363134
rect 354606 362898 385090 363134
rect 385326 362898 415810 363134
rect 416046 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 586890 363134
rect -2966 362866 586890 362898
rect -8726 356614 592650 356646
rect -8726 356378 -8694 356614
rect -8458 356378 -8374 356614
rect -8138 356378 30986 356614
rect 31222 356378 31306 356614
rect 31542 356378 66986 356614
rect 67222 356378 67306 356614
rect 67542 356378 102986 356614
rect 103222 356378 103306 356614
rect 103542 356378 138986 356614
rect 139222 356378 139306 356614
rect 139542 356378 426986 356614
rect 427222 356378 427306 356614
rect 427542 356378 462986 356614
rect 463222 356378 463306 356614
rect 463542 356378 498986 356614
rect 499222 356378 499306 356614
rect 499542 356378 534986 356614
rect 535222 356378 535306 356614
rect 535542 356378 570986 356614
rect 571222 356378 571306 356614
rect 571542 356378 592062 356614
rect 592298 356378 592382 356614
rect 592618 356378 592650 356614
rect -8726 356294 592650 356378
rect -8726 356058 -8694 356294
rect -8458 356058 -8374 356294
rect -8138 356058 30986 356294
rect 31222 356058 31306 356294
rect 31542 356058 66986 356294
rect 67222 356058 67306 356294
rect 67542 356058 102986 356294
rect 103222 356058 103306 356294
rect 103542 356058 138986 356294
rect 139222 356058 139306 356294
rect 139542 356058 426986 356294
rect 427222 356058 427306 356294
rect 427542 356058 462986 356294
rect 463222 356058 463306 356294
rect 463542 356058 498986 356294
rect 499222 356058 499306 356294
rect 499542 356058 534986 356294
rect 535222 356058 535306 356294
rect 535542 356058 570986 356294
rect 571222 356058 571306 356294
rect 571542 356058 592062 356294
rect 592298 356058 592382 356294
rect 592618 356058 592650 356294
rect -8726 356026 592650 356058
rect -6806 352894 590730 352926
rect -6806 352658 -6774 352894
rect -6538 352658 -6454 352894
rect -6218 352658 27266 352894
rect 27502 352658 27586 352894
rect 27822 352658 63266 352894
rect 63502 352658 63586 352894
rect 63822 352658 99266 352894
rect 99502 352658 99586 352894
rect 99822 352658 135266 352894
rect 135502 352658 135586 352894
rect 135822 352658 423266 352894
rect 423502 352658 423586 352894
rect 423822 352658 459266 352894
rect 459502 352658 459586 352894
rect 459822 352658 495266 352894
rect 495502 352658 495586 352894
rect 495822 352658 531266 352894
rect 531502 352658 531586 352894
rect 531822 352658 567266 352894
rect 567502 352658 567586 352894
rect 567822 352658 590142 352894
rect 590378 352658 590462 352894
rect 590698 352658 590730 352894
rect -6806 352574 590730 352658
rect -6806 352338 -6774 352574
rect -6538 352338 -6454 352574
rect -6218 352338 27266 352574
rect 27502 352338 27586 352574
rect 27822 352338 63266 352574
rect 63502 352338 63586 352574
rect 63822 352338 99266 352574
rect 99502 352338 99586 352574
rect 99822 352338 135266 352574
rect 135502 352338 135586 352574
rect 135822 352338 423266 352574
rect 423502 352338 423586 352574
rect 423822 352338 459266 352574
rect 459502 352338 459586 352574
rect 459822 352338 495266 352574
rect 495502 352338 495586 352574
rect 495822 352338 531266 352574
rect 531502 352338 531586 352574
rect 531822 352338 567266 352574
rect 567502 352338 567586 352574
rect 567822 352338 590142 352574
rect 590378 352338 590462 352574
rect 590698 352338 590730 352574
rect -6806 352306 590730 352338
rect -4886 349174 588810 349206
rect -4886 348938 -4854 349174
rect -4618 348938 -4534 349174
rect -4298 348938 23546 349174
rect 23782 348938 23866 349174
rect 24102 348938 59546 349174
rect 59782 348938 59866 349174
rect 60102 348938 95546 349174
rect 95782 348938 95866 349174
rect 96102 348938 131546 349174
rect 131782 348938 131866 349174
rect 132102 348938 455546 349174
rect 455782 348938 455866 349174
rect 456102 348938 491546 349174
rect 491782 348938 491866 349174
rect 492102 348938 527546 349174
rect 527782 348938 527866 349174
rect 528102 348938 563546 349174
rect 563782 348938 563866 349174
rect 564102 348938 588222 349174
rect 588458 348938 588542 349174
rect 588778 348938 588810 349174
rect -4886 348854 588810 348938
rect -4886 348618 -4854 348854
rect -4618 348618 -4534 348854
rect -4298 348618 23546 348854
rect 23782 348618 23866 348854
rect 24102 348618 59546 348854
rect 59782 348618 59866 348854
rect 60102 348618 95546 348854
rect 95782 348618 95866 348854
rect 96102 348618 131546 348854
rect 131782 348618 131866 348854
rect 132102 348618 455546 348854
rect 455782 348618 455866 348854
rect 456102 348618 491546 348854
rect 491782 348618 491866 348854
rect 492102 348618 527546 348854
rect 527782 348618 527866 348854
rect 528102 348618 563546 348854
rect 563782 348618 563866 348854
rect 564102 348618 588222 348854
rect 588458 348618 588542 348854
rect 588778 348618 588810 348854
rect -4886 348586 588810 348618
rect -2966 345454 586890 345486
rect -2966 345218 -2934 345454
rect -2698 345218 -2614 345454
rect -2378 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 91826 345454
rect 92062 345218 92146 345454
rect 92382 345218 127826 345454
rect 128062 345218 128146 345454
rect 128382 345218 185410 345454
rect 185646 345218 216130 345454
rect 216366 345218 246850 345454
rect 247086 345218 277570 345454
rect 277806 345218 308290 345454
rect 308526 345218 339010 345454
rect 339246 345218 369730 345454
rect 369966 345218 400450 345454
rect 400686 345218 451826 345454
rect 452062 345218 452146 345454
rect 452382 345218 487826 345454
rect 488062 345218 488146 345454
rect 488382 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 586302 345454
rect 586538 345218 586622 345454
rect 586858 345218 586890 345454
rect -2966 345134 586890 345218
rect -2966 344898 -2934 345134
rect -2698 344898 -2614 345134
rect -2378 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 91826 345134
rect 92062 344898 92146 345134
rect 92382 344898 127826 345134
rect 128062 344898 128146 345134
rect 128382 344898 185410 345134
rect 185646 344898 216130 345134
rect 216366 344898 246850 345134
rect 247086 344898 277570 345134
rect 277806 344898 308290 345134
rect 308526 344898 339010 345134
rect 339246 344898 369730 345134
rect 369966 344898 400450 345134
rect 400686 344898 451826 345134
rect 452062 344898 452146 345134
rect 452382 344898 487826 345134
rect 488062 344898 488146 345134
rect 488382 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 586302 345134
rect 586538 344898 586622 345134
rect 586858 344898 586890 345134
rect -2966 344866 586890 344898
rect -8726 338614 592650 338646
rect -8726 338378 -7734 338614
rect -7498 338378 -7414 338614
rect -7178 338378 12986 338614
rect 13222 338378 13306 338614
rect 13542 338378 48986 338614
rect 49222 338378 49306 338614
rect 49542 338378 84986 338614
rect 85222 338378 85306 338614
rect 85542 338378 120986 338614
rect 121222 338378 121306 338614
rect 121542 338378 156986 338614
rect 157222 338378 157306 338614
rect 157542 338378 444986 338614
rect 445222 338378 445306 338614
rect 445542 338378 480986 338614
rect 481222 338378 481306 338614
rect 481542 338378 516986 338614
rect 517222 338378 517306 338614
rect 517542 338378 552986 338614
rect 553222 338378 553306 338614
rect 553542 338378 591102 338614
rect 591338 338378 591422 338614
rect 591658 338378 592650 338614
rect -8726 338294 592650 338378
rect -8726 338058 -7734 338294
rect -7498 338058 -7414 338294
rect -7178 338058 12986 338294
rect 13222 338058 13306 338294
rect 13542 338058 48986 338294
rect 49222 338058 49306 338294
rect 49542 338058 84986 338294
rect 85222 338058 85306 338294
rect 85542 338058 120986 338294
rect 121222 338058 121306 338294
rect 121542 338058 156986 338294
rect 157222 338058 157306 338294
rect 157542 338058 444986 338294
rect 445222 338058 445306 338294
rect 445542 338058 480986 338294
rect 481222 338058 481306 338294
rect 481542 338058 516986 338294
rect 517222 338058 517306 338294
rect 517542 338058 552986 338294
rect 553222 338058 553306 338294
rect 553542 338058 591102 338294
rect 591338 338058 591422 338294
rect 591658 338058 592650 338294
rect -8726 338026 592650 338058
rect -6806 334894 590730 334926
rect -6806 334658 -5814 334894
rect -5578 334658 -5494 334894
rect -5258 334658 9266 334894
rect 9502 334658 9586 334894
rect 9822 334658 45266 334894
rect 45502 334658 45586 334894
rect 45822 334658 81266 334894
rect 81502 334658 81586 334894
rect 81822 334658 117266 334894
rect 117502 334658 117586 334894
rect 117822 334658 153266 334894
rect 153502 334658 153586 334894
rect 153822 334658 441266 334894
rect 441502 334658 441586 334894
rect 441822 334658 477266 334894
rect 477502 334658 477586 334894
rect 477822 334658 513266 334894
rect 513502 334658 513586 334894
rect 513822 334658 549266 334894
rect 549502 334658 549586 334894
rect 549822 334658 589182 334894
rect 589418 334658 589502 334894
rect 589738 334658 590730 334894
rect -6806 334574 590730 334658
rect -6806 334338 -5814 334574
rect -5578 334338 -5494 334574
rect -5258 334338 9266 334574
rect 9502 334338 9586 334574
rect 9822 334338 45266 334574
rect 45502 334338 45586 334574
rect 45822 334338 81266 334574
rect 81502 334338 81586 334574
rect 81822 334338 117266 334574
rect 117502 334338 117586 334574
rect 117822 334338 153266 334574
rect 153502 334338 153586 334574
rect 153822 334338 441266 334574
rect 441502 334338 441586 334574
rect 441822 334338 477266 334574
rect 477502 334338 477586 334574
rect 477822 334338 513266 334574
rect 513502 334338 513586 334574
rect 513822 334338 549266 334574
rect 549502 334338 549586 334574
rect 549822 334338 589182 334574
rect 589418 334338 589502 334574
rect 589738 334338 590730 334574
rect -6806 334306 590730 334338
rect -4886 331174 588810 331206
rect -4886 330938 -3894 331174
rect -3658 330938 -3574 331174
rect -3338 330938 5546 331174
rect 5782 330938 5866 331174
rect 6102 330938 41546 331174
rect 41782 330938 41866 331174
rect 42102 330938 77546 331174
rect 77782 330938 77866 331174
rect 78102 330938 113546 331174
rect 113782 330938 113866 331174
rect 114102 330938 149546 331174
rect 149782 330938 149866 331174
rect 150102 330938 437546 331174
rect 437782 330938 437866 331174
rect 438102 330938 473546 331174
rect 473782 330938 473866 331174
rect 474102 330938 509546 331174
rect 509782 330938 509866 331174
rect 510102 330938 545546 331174
rect 545782 330938 545866 331174
rect 546102 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 587262 331174
rect 587498 330938 587582 331174
rect 587818 330938 588810 331174
rect -4886 330854 588810 330938
rect -4886 330618 -3894 330854
rect -3658 330618 -3574 330854
rect -3338 330618 5546 330854
rect 5782 330618 5866 330854
rect 6102 330618 41546 330854
rect 41782 330618 41866 330854
rect 42102 330618 77546 330854
rect 77782 330618 77866 330854
rect 78102 330618 113546 330854
rect 113782 330618 113866 330854
rect 114102 330618 149546 330854
rect 149782 330618 149866 330854
rect 150102 330618 437546 330854
rect 437782 330618 437866 330854
rect 438102 330618 473546 330854
rect 473782 330618 473866 330854
rect 474102 330618 509546 330854
rect 509782 330618 509866 330854
rect 510102 330618 545546 330854
rect 545782 330618 545866 330854
rect 546102 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 587262 330854
rect 587498 330618 587582 330854
rect 587818 330618 588810 330854
rect -4886 330586 588810 330618
rect -2966 327454 586890 327486
rect -2966 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 73826 327454
rect 74062 327218 74146 327454
rect 74382 327218 109826 327454
rect 110062 327218 110146 327454
rect 110382 327218 145826 327454
rect 146062 327218 146146 327454
rect 146382 327218 170050 327454
rect 170286 327218 200770 327454
rect 201006 327218 231490 327454
rect 231726 327218 262210 327454
rect 262446 327218 292930 327454
rect 293166 327218 323650 327454
rect 323886 327218 354370 327454
rect 354606 327218 385090 327454
rect 385326 327218 415810 327454
rect 416046 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 586890 327454
rect -2966 327134 586890 327218
rect -2966 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 73826 327134
rect 74062 326898 74146 327134
rect 74382 326898 109826 327134
rect 110062 326898 110146 327134
rect 110382 326898 145826 327134
rect 146062 326898 146146 327134
rect 146382 326898 170050 327134
rect 170286 326898 200770 327134
rect 201006 326898 231490 327134
rect 231726 326898 262210 327134
rect 262446 326898 292930 327134
rect 293166 326898 323650 327134
rect 323886 326898 354370 327134
rect 354606 326898 385090 327134
rect 385326 326898 415810 327134
rect 416046 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 586890 327134
rect -2966 326866 586890 326898
rect -8726 320614 592650 320646
rect -8726 320378 -8694 320614
rect -8458 320378 -8374 320614
rect -8138 320378 30986 320614
rect 31222 320378 31306 320614
rect 31542 320378 66986 320614
rect 67222 320378 67306 320614
rect 67542 320378 102986 320614
rect 103222 320378 103306 320614
rect 103542 320378 138986 320614
rect 139222 320378 139306 320614
rect 139542 320378 426986 320614
rect 427222 320378 427306 320614
rect 427542 320378 462986 320614
rect 463222 320378 463306 320614
rect 463542 320378 498986 320614
rect 499222 320378 499306 320614
rect 499542 320378 534986 320614
rect 535222 320378 535306 320614
rect 535542 320378 570986 320614
rect 571222 320378 571306 320614
rect 571542 320378 592062 320614
rect 592298 320378 592382 320614
rect 592618 320378 592650 320614
rect -8726 320294 592650 320378
rect -8726 320058 -8694 320294
rect -8458 320058 -8374 320294
rect -8138 320058 30986 320294
rect 31222 320058 31306 320294
rect 31542 320058 66986 320294
rect 67222 320058 67306 320294
rect 67542 320058 102986 320294
rect 103222 320058 103306 320294
rect 103542 320058 138986 320294
rect 139222 320058 139306 320294
rect 139542 320058 426986 320294
rect 427222 320058 427306 320294
rect 427542 320058 462986 320294
rect 463222 320058 463306 320294
rect 463542 320058 498986 320294
rect 499222 320058 499306 320294
rect 499542 320058 534986 320294
rect 535222 320058 535306 320294
rect 535542 320058 570986 320294
rect 571222 320058 571306 320294
rect 571542 320058 592062 320294
rect 592298 320058 592382 320294
rect 592618 320058 592650 320294
rect -8726 320026 592650 320058
rect -6806 316894 590730 316926
rect -6806 316658 -6774 316894
rect -6538 316658 -6454 316894
rect -6218 316658 27266 316894
rect 27502 316658 27586 316894
rect 27822 316658 63266 316894
rect 63502 316658 63586 316894
rect 63822 316658 99266 316894
rect 99502 316658 99586 316894
rect 99822 316658 135266 316894
rect 135502 316658 135586 316894
rect 135822 316658 423266 316894
rect 423502 316658 423586 316894
rect 423822 316658 459266 316894
rect 459502 316658 459586 316894
rect 459822 316658 495266 316894
rect 495502 316658 495586 316894
rect 495822 316658 531266 316894
rect 531502 316658 531586 316894
rect 531822 316658 567266 316894
rect 567502 316658 567586 316894
rect 567822 316658 590142 316894
rect 590378 316658 590462 316894
rect 590698 316658 590730 316894
rect -6806 316574 590730 316658
rect -6806 316338 -6774 316574
rect -6538 316338 -6454 316574
rect -6218 316338 27266 316574
rect 27502 316338 27586 316574
rect 27822 316338 63266 316574
rect 63502 316338 63586 316574
rect 63822 316338 99266 316574
rect 99502 316338 99586 316574
rect 99822 316338 135266 316574
rect 135502 316338 135586 316574
rect 135822 316338 423266 316574
rect 423502 316338 423586 316574
rect 423822 316338 459266 316574
rect 459502 316338 459586 316574
rect 459822 316338 495266 316574
rect 495502 316338 495586 316574
rect 495822 316338 531266 316574
rect 531502 316338 531586 316574
rect 531822 316338 567266 316574
rect 567502 316338 567586 316574
rect 567822 316338 590142 316574
rect 590378 316338 590462 316574
rect 590698 316338 590730 316574
rect -6806 316306 590730 316338
rect -4886 313174 588810 313206
rect -4886 312938 -4854 313174
rect -4618 312938 -4534 313174
rect -4298 312938 23546 313174
rect 23782 312938 23866 313174
rect 24102 312938 59546 313174
rect 59782 312938 59866 313174
rect 60102 312938 95546 313174
rect 95782 312938 95866 313174
rect 96102 312938 131546 313174
rect 131782 312938 131866 313174
rect 132102 312938 455546 313174
rect 455782 312938 455866 313174
rect 456102 312938 491546 313174
rect 491782 312938 491866 313174
rect 492102 312938 527546 313174
rect 527782 312938 527866 313174
rect 528102 312938 563546 313174
rect 563782 312938 563866 313174
rect 564102 312938 588222 313174
rect 588458 312938 588542 313174
rect 588778 312938 588810 313174
rect -4886 312854 588810 312938
rect -4886 312618 -4854 312854
rect -4618 312618 -4534 312854
rect -4298 312618 23546 312854
rect 23782 312618 23866 312854
rect 24102 312618 59546 312854
rect 59782 312618 59866 312854
rect 60102 312618 95546 312854
rect 95782 312618 95866 312854
rect 96102 312618 131546 312854
rect 131782 312618 131866 312854
rect 132102 312618 455546 312854
rect 455782 312618 455866 312854
rect 456102 312618 491546 312854
rect 491782 312618 491866 312854
rect 492102 312618 527546 312854
rect 527782 312618 527866 312854
rect 528102 312618 563546 312854
rect 563782 312618 563866 312854
rect 564102 312618 588222 312854
rect 588458 312618 588542 312854
rect 588778 312618 588810 312854
rect -4886 312586 588810 312618
rect -2966 309454 586890 309486
rect -2966 309218 -2934 309454
rect -2698 309218 -2614 309454
rect -2378 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 91826 309454
rect 92062 309218 92146 309454
rect 92382 309218 127826 309454
rect 128062 309218 128146 309454
rect 128382 309218 185410 309454
rect 185646 309218 216130 309454
rect 216366 309218 246850 309454
rect 247086 309218 277570 309454
rect 277806 309218 308290 309454
rect 308526 309218 339010 309454
rect 339246 309218 369730 309454
rect 369966 309218 400450 309454
rect 400686 309218 451826 309454
rect 452062 309218 452146 309454
rect 452382 309218 487826 309454
rect 488062 309218 488146 309454
rect 488382 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 586302 309454
rect 586538 309218 586622 309454
rect 586858 309218 586890 309454
rect -2966 309134 586890 309218
rect -2966 308898 -2934 309134
rect -2698 308898 -2614 309134
rect -2378 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 91826 309134
rect 92062 308898 92146 309134
rect 92382 308898 127826 309134
rect 128062 308898 128146 309134
rect 128382 308898 185410 309134
rect 185646 308898 216130 309134
rect 216366 308898 246850 309134
rect 247086 308898 277570 309134
rect 277806 308898 308290 309134
rect 308526 308898 339010 309134
rect 339246 308898 369730 309134
rect 369966 308898 400450 309134
rect 400686 308898 451826 309134
rect 452062 308898 452146 309134
rect 452382 308898 487826 309134
rect 488062 308898 488146 309134
rect 488382 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 586302 309134
rect 586538 308898 586622 309134
rect 586858 308898 586890 309134
rect -2966 308866 586890 308898
rect -8726 302614 592650 302646
rect -8726 302378 -7734 302614
rect -7498 302378 -7414 302614
rect -7178 302378 12986 302614
rect 13222 302378 13306 302614
rect 13542 302378 48986 302614
rect 49222 302378 49306 302614
rect 49542 302378 84986 302614
rect 85222 302378 85306 302614
rect 85542 302378 120986 302614
rect 121222 302378 121306 302614
rect 121542 302378 156986 302614
rect 157222 302378 157306 302614
rect 157542 302378 444986 302614
rect 445222 302378 445306 302614
rect 445542 302378 480986 302614
rect 481222 302378 481306 302614
rect 481542 302378 516986 302614
rect 517222 302378 517306 302614
rect 517542 302378 552986 302614
rect 553222 302378 553306 302614
rect 553542 302378 591102 302614
rect 591338 302378 591422 302614
rect 591658 302378 592650 302614
rect -8726 302294 592650 302378
rect -8726 302058 -7734 302294
rect -7498 302058 -7414 302294
rect -7178 302058 12986 302294
rect 13222 302058 13306 302294
rect 13542 302058 48986 302294
rect 49222 302058 49306 302294
rect 49542 302058 84986 302294
rect 85222 302058 85306 302294
rect 85542 302058 120986 302294
rect 121222 302058 121306 302294
rect 121542 302058 156986 302294
rect 157222 302058 157306 302294
rect 157542 302058 444986 302294
rect 445222 302058 445306 302294
rect 445542 302058 480986 302294
rect 481222 302058 481306 302294
rect 481542 302058 516986 302294
rect 517222 302058 517306 302294
rect 517542 302058 552986 302294
rect 553222 302058 553306 302294
rect 553542 302058 591102 302294
rect 591338 302058 591422 302294
rect 591658 302058 592650 302294
rect -8726 302026 592650 302058
rect -6806 298894 590730 298926
rect -6806 298658 -5814 298894
rect -5578 298658 -5494 298894
rect -5258 298658 9266 298894
rect 9502 298658 9586 298894
rect 9822 298658 45266 298894
rect 45502 298658 45586 298894
rect 45822 298658 81266 298894
rect 81502 298658 81586 298894
rect 81822 298658 117266 298894
rect 117502 298658 117586 298894
rect 117822 298658 153266 298894
rect 153502 298658 153586 298894
rect 153822 298658 441266 298894
rect 441502 298658 441586 298894
rect 441822 298658 477266 298894
rect 477502 298658 477586 298894
rect 477822 298658 513266 298894
rect 513502 298658 513586 298894
rect 513822 298658 549266 298894
rect 549502 298658 549586 298894
rect 549822 298658 589182 298894
rect 589418 298658 589502 298894
rect 589738 298658 590730 298894
rect -6806 298574 590730 298658
rect -6806 298338 -5814 298574
rect -5578 298338 -5494 298574
rect -5258 298338 9266 298574
rect 9502 298338 9586 298574
rect 9822 298338 45266 298574
rect 45502 298338 45586 298574
rect 45822 298338 81266 298574
rect 81502 298338 81586 298574
rect 81822 298338 117266 298574
rect 117502 298338 117586 298574
rect 117822 298338 153266 298574
rect 153502 298338 153586 298574
rect 153822 298338 441266 298574
rect 441502 298338 441586 298574
rect 441822 298338 477266 298574
rect 477502 298338 477586 298574
rect 477822 298338 513266 298574
rect 513502 298338 513586 298574
rect 513822 298338 549266 298574
rect 549502 298338 549586 298574
rect 549822 298338 589182 298574
rect 589418 298338 589502 298574
rect 589738 298338 590730 298574
rect -6806 298306 590730 298338
rect -4886 295174 588810 295206
rect -4886 294938 -3894 295174
rect -3658 294938 -3574 295174
rect -3338 294938 5546 295174
rect 5782 294938 5866 295174
rect 6102 294938 41546 295174
rect 41782 294938 41866 295174
rect 42102 294938 77546 295174
rect 77782 294938 77866 295174
rect 78102 294938 113546 295174
rect 113782 294938 113866 295174
rect 114102 294938 149546 295174
rect 149782 294938 149866 295174
rect 150102 294938 437546 295174
rect 437782 294938 437866 295174
rect 438102 294938 473546 295174
rect 473782 294938 473866 295174
rect 474102 294938 509546 295174
rect 509782 294938 509866 295174
rect 510102 294938 545546 295174
rect 545782 294938 545866 295174
rect 546102 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 587262 295174
rect 587498 294938 587582 295174
rect 587818 294938 588810 295174
rect -4886 294854 588810 294938
rect -4886 294618 -3894 294854
rect -3658 294618 -3574 294854
rect -3338 294618 5546 294854
rect 5782 294618 5866 294854
rect 6102 294618 41546 294854
rect 41782 294618 41866 294854
rect 42102 294618 77546 294854
rect 77782 294618 77866 294854
rect 78102 294618 113546 294854
rect 113782 294618 113866 294854
rect 114102 294618 149546 294854
rect 149782 294618 149866 294854
rect 150102 294618 437546 294854
rect 437782 294618 437866 294854
rect 438102 294618 473546 294854
rect 473782 294618 473866 294854
rect 474102 294618 509546 294854
rect 509782 294618 509866 294854
rect 510102 294618 545546 294854
rect 545782 294618 545866 294854
rect 546102 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 587262 294854
rect 587498 294618 587582 294854
rect 587818 294618 588810 294854
rect -4886 294586 588810 294618
rect -2966 291454 586890 291486
rect -2966 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 73826 291454
rect 74062 291218 74146 291454
rect 74382 291218 109826 291454
rect 110062 291218 110146 291454
rect 110382 291218 145826 291454
rect 146062 291218 146146 291454
rect 146382 291218 170050 291454
rect 170286 291218 200770 291454
rect 201006 291218 231490 291454
rect 231726 291218 262210 291454
rect 262446 291218 292930 291454
rect 293166 291218 323650 291454
rect 323886 291218 354370 291454
rect 354606 291218 385090 291454
rect 385326 291218 415810 291454
rect 416046 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 586890 291454
rect -2966 291134 586890 291218
rect -2966 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 73826 291134
rect 74062 290898 74146 291134
rect 74382 290898 109826 291134
rect 110062 290898 110146 291134
rect 110382 290898 145826 291134
rect 146062 290898 146146 291134
rect 146382 290898 170050 291134
rect 170286 290898 200770 291134
rect 201006 290898 231490 291134
rect 231726 290898 262210 291134
rect 262446 290898 292930 291134
rect 293166 290898 323650 291134
rect 323886 290898 354370 291134
rect 354606 290898 385090 291134
rect 385326 290898 415810 291134
rect 416046 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 586890 291134
rect -2966 290866 586890 290898
rect -8726 284614 592650 284646
rect -8726 284378 -8694 284614
rect -8458 284378 -8374 284614
rect -8138 284378 30986 284614
rect 31222 284378 31306 284614
rect 31542 284378 66986 284614
rect 67222 284378 67306 284614
rect 67542 284378 102986 284614
rect 103222 284378 103306 284614
rect 103542 284378 138986 284614
rect 139222 284378 139306 284614
rect 139542 284378 426986 284614
rect 427222 284378 427306 284614
rect 427542 284378 462986 284614
rect 463222 284378 463306 284614
rect 463542 284378 498986 284614
rect 499222 284378 499306 284614
rect 499542 284378 534986 284614
rect 535222 284378 535306 284614
rect 535542 284378 570986 284614
rect 571222 284378 571306 284614
rect 571542 284378 592062 284614
rect 592298 284378 592382 284614
rect 592618 284378 592650 284614
rect -8726 284294 592650 284378
rect -8726 284058 -8694 284294
rect -8458 284058 -8374 284294
rect -8138 284058 30986 284294
rect 31222 284058 31306 284294
rect 31542 284058 66986 284294
rect 67222 284058 67306 284294
rect 67542 284058 102986 284294
rect 103222 284058 103306 284294
rect 103542 284058 138986 284294
rect 139222 284058 139306 284294
rect 139542 284058 426986 284294
rect 427222 284058 427306 284294
rect 427542 284058 462986 284294
rect 463222 284058 463306 284294
rect 463542 284058 498986 284294
rect 499222 284058 499306 284294
rect 499542 284058 534986 284294
rect 535222 284058 535306 284294
rect 535542 284058 570986 284294
rect 571222 284058 571306 284294
rect 571542 284058 592062 284294
rect 592298 284058 592382 284294
rect 592618 284058 592650 284294
rect -8726 284026 592650 284058
rect -6806 280894 590730 280926
rect -6806 280658 -6774 280894
rect -6538 280658 -6454 280894
rect -6218 280658 27266 280894
rect 27502 280658 27586 280894
rect 27822 280658 63266 280894
rect 63502 280658 63586 280894
rect 63822 280658 99266 280894
rect 99502 280658 99586 280894
rect 99822 280658 135266 280894
rect 135502 280658 135586 280894
rect 135822 280658 423266 280894
rect 423502 280658 423586 280894
rect 423822 280658 459266 280894
rect 459502 280658 459586 280894
rect 459822 280658 495266 280894
rect 495502 280658 495586 280894
rect 495822 280658 531266 280894
rect 531502 280658 531586 280894
rect 531822 280658 567266 280894
rect 567502 280658 567586 280894
rect 567822 280658 590142 280894
rect 590378 280658 590462 280894
rect 590698 280658 590730 280894
rect -6806 280574 590730 280658
rect -6806 280338 -6774 280574
rect -6538 280338 -6454 280574
rect -6218 280338 27266 280574
rect 27502 280338 27586 280574
rect 27822 280338 63266 280574
rect 63502 280338 63586 280574
rect 63822 280338 99266 280574
rect 99502 280338 99586 280574
rect 99822 280338 135266 280574
rect 135502 280338 135586 280574
rect 135822 280338 423266 280574
rect 423502 280338 423586 280574
rect 423822 280338 459266 280574
rect 459502 280338 459586 280574
rect 459822 280338 495266 280574
rect 495502 280338 495586 280574
rect 495822 280338 531266 280574
rect 531502 280338 531586 280574
rect 531822 280338 567266 280574
rect 567502 280338 567586 280574
rect 567822 280338 590142 280574
rect 590378 280338 590462 280574
rect 590698 280338 590730 280574
rect -6806 280306 590730 280338
rect -4886 277174 588810 277206
rect -4886 276938 -4854 277174
rect -4618 276938 -4534 277174
rect -4298 276938 23546 277174
rect 23782 276938 23866 277174
rect 24102 276938 59546 277174
rect 59782 276938 59866 277174
rect 60102 276938 95546 277174
rect 95782 276938 95866 277174
rect 96102 276938 131546 277174
rect 131782 276938 131866 277174
rect 132102 276938 455546 277174
rect 455782 276938 455866 277174
rect 456102 276938 491546 277174
rect 491782 276938 491866 277174
rect 492102 276938 527546 277174
rect 527782 276938 527866 277174
rect 528102 276938 563546 277174
rect 563782 276938 563866 277174
rect 564102 276938 588222 277174
rect 588458 276938 588542 277174
rect 588778 276938 588810 277174
rect -4886 276854 588810 276938
rect -4886 276618 -4854 276854
rect -4618 276618 -4534 276854
rect -4298 276618 23546 276854
rect 23782 276618 23866 276854
rect 24102 276618 59546 276854
rect 59782 276618 59866 276854
rect 60102 276618 95546 276854
rect 95782 276618 95866 276854
rect 96102 276618 131546 276854
rect 131782 276618 131866 276854
rect 132102 276618 455546 276854
rect 455782 276618 455866 276854
rect 456102 276618 491546 276854
rect 491782 276618 491866 276854
rect 492102 276618 527546 276854
rect 527782 276618 527866 276854
rect 528102 276618 563546 276854
rect 563782 276618 563866 276854
rect 564102 276618 588222 276854
rect 588458 276618 588542 276854
rect 588778 276618 588810 276854
rect -4886 276586 588810 276618
rect -2966 273454 586890 273486
rect -2966 273218 -2934 273454
rect -2698 273218 -2614 273454
rect -2378 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 91826 273454
rect 92062 273218 92146 273454
rect 92382 273218 127826 273454
rect 128062 273218 128146 273454
rect 128382 273218 185410 273454
rect 185646 273218 216130 273454
rect 216366 273218 246850 273454
rect 247086 273218 277570 273454
rect 277806 273218 308290 273454
rect 308526 273218 339010 273454
rect 339246 273218 369730 273454
rect 369966 273218 400450 273454
rect 400686 273218 451826 273454
rect 452062 273218 452146 273454
rect 452382 273218 487826 273454
rect 488062 273218 488146 273454
rect 488382 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 586302 273454
rect 586538 273218 586622 273454
rect 586858 273218 586890 273454
rect -2966 273134 586890 273218
rect -2966 272898 -2934 273134
rect -2698 272898 -2614 273134
rect -2378 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 91826 273134
rect 92062 272898 92146 273134
rect 92382 272898 127826 273134
rect 128062 272898 128146 273134
rect 128382 272898 185410 273134
rect 185646 272898 216130 273134
rect 216366 272898 246850 273134
rect 247086 272898 277570 273134
rect 277806 272898 308290 273134
rect 308526 272898 339010 273134
rect 339246 272898 369730 273134
rect 369966 272898 400450 273134
rect 400686 272898 451826 273134
rect 452062 272898 452146 273134
rect 452382 272898 487826 273134
rect 488062 272898 488146 273134
rect 488382 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 586302 273134
rect 586538 272898 586622 273134
rect 586858 272898 586890 273134
rect -2966 272866 586890 272898
rect -8726 266614 592650 266646
rect -8726 266378 -7734 266614
rect -7498 266378 -7414 266614
rect -7178 266378 12986 266614
rect 13222 266378 13306 266614
rect 13542 266378 48986 266614
rect 49222 266378 49306 266614
rect 49542 266378 84986 266614
rect 85222 266378 85306 266614
rect 85542 266378 120986 266614
rect 121222 266378 121306 266614
rect 121542 266378 156986 266614
rect 157222 266378 157306 266614
rect 157542 266378 444986 266614
rect 445222 266378 445306 266614
rect 445542 266378 480986 266614
rect 481222 266378 481306 266614
rect 481542 266378 516986 266614
rect 517222 266378 517306 266614
rect 517542 266378 552986 266614
rect 553222 266378 553306 266614
rect 553542 266378 591102 266614
rect 591338 266378 591422 266614
rect 591658 266378 592650 266614
rect -8726 266294 592650 266378
rect -8726 266058 -7734 266294
rect -7498 266058 -7414 266294
rect -7178 266058 12986 266294
rect 13222 266058 13306 266294
rect 13542 266058 48986 266294
rect 49222 266058 49306 266294
rect 49542 266058 84986 266294
rect 85222 266058 85306 266294
rect 85542 266058 120986 266294
rect 121222 266058 121306 266294
rect 121542 266058 156986 266294
rect 157222 266058 157306 266294
rect 157542 266058 444986 266294
rect 445222 266058 445306 266294
rect 445542 266058 480986 266294
rect 481222 266058 481306 266294
rect 481542 266058 516986 266294
rect 517222 266058 517306 266294
rect 517542 266058 552986 266294
rect 553222 266058 553306 266294
rect 553542 266058 591102 266294
rect 591338 266058 591422 266294
rect 591658 266058 592650 266294
rect -8726 266026 592650 266058
rect -6806 262894 590730 262926
rect -6806 262658 -5814 262894
rect -5578 262658 -5494 262894
rect -5258 262658 9266 262894
rect 9502 262658 9586 262894
rect 9822 262658 45266 262894
rect 45502 262658 45586 262894
rect 45822 262658 81266 262894
rect 81502 262658 81586 262894
rect 81822 262658 117266 262894
rect 117502 262658 117586 262894
rect 117822 262658 153266 262894
rect 153502 262658 153586 262894
rect 153822 262658 441266 262894
rect 441502 262658 441586 262894
rect 441822 262658 477266 262894
rect 477502 262658 477586 262894
rect 477822 262658 513266 262894
rect 513502 262658 513586 262894
rect 513822 262658 549266 262894
rect 549502 262658 549586 262894
rect 549822 262658 589182 262894
rect 589418 262658 589502 262894
rect 589738 262658 590730 262894
rect -6806 262574 590730 262658
rect -6806 262338 -5814 262574
rect -5578 262338 -5494 262574
rect -5258 262338 9266 262574
rect 9502 262338 9586 262574
rect 9822 262338 45266 262574
rect 45502 262338 45586 262574
rect 45822 262338 81266 262574
rect 81502 262338 81586 262574
rect 81822 262338 117266 262574
rect 117502 262338 117586 262574
rect 117822 262338 153266 262574
rect 153502 262338 153586 262574
rect 153822 262338 441266 262574
rect 441502 262338 441586 262574
rect 441822 262338 477266 262574
rect 477502 262338 477586 262574
rect 477822 262338 513266 262574
rect 513502 262338 513586 262574
rect 513822 262338 549266 262574
rect 549502 262338 549586 262574
rect 549822 262338 589182 262574
rect 589418 262338 589502 262574
rect 589738 262338 590730 262574
rect -6806 262306 590730 262338
rect -4886 259174 588810 259206
rect -4886 258938 -3894 259174
rect -3658 258938 -3574 259174
rect -3338 258938 5546 259174
rect 5782 258938 5866 259174
rect 6102 258938 41546 259174
rect 41782 258938 41866 259174
rect 42102 258938 77546 259174
rect 77782 258938 77866 259174
rect 78102 258938 113546 259174
rect 113782 258938 113866 259174
rect 114102 258938 149546 259174
rect 149782 258938 149866 259174
rect 150102 258938 437546 259174
rect 437782 258938 437866 259174
rect 438102 258938 473546 259174
rect 473782 258938 473866 259174
rect 474102 258938 509546 259174
rect 509782 258938 509866 259174
rect 510102 258938 545546 259174
rect 545782 258938 545866 259174
rect 546102 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 587262 259174
rect 587498 258938 587582 259174
rect 587818 258938 588810 259174
rect -4886 258854 588810 258938
rect -4886 258618 -3894 258854
rect -3658 258618 -3574 258854
rect -3338 258618 5546 258854
rect 5782 258618 5866 258854
rect 6102 258618 41546 258854
rect 41782 258618 41866 258854
rect 42102 258618 77546 258854
rect 77782 258618 77866 258854
rect 78102 258618 113546 258854
rect 113782 258618 113866 258854
rect 114102 258618 149546 258854
rect 149782 258618 149866 258854
rect 150102 258618 437546 258854
rect 437782 258618 437866 258854
rect 438102 258618 473546 258854
rect 473782 258618 473866 258854
rect 474102 258618 509546 258854
rect 509782 258618 509866 258854
rect 510102 258618 545546 258854
rect 545782 258618 545866 258854
rect 546102 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 587262 258854
rect 587498 258618 587582 258854
rect 587818 258618 588810 258854
rect -4886 258586 588810 258618
rect -2966 255454 586890 255486
rect -2966 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 73826 255454
rect 74062 255218 74146 255454
rect 74382 255218 109826 255454
rect 110062 255218 110146 255454
rect 110382 255218 145826 255454
rect 146062 255218 146146 255454
rect 146382 255218 170050 255454
rect 170286 255218 200770 255454
rect 201006 255218 231490 255454
rect 231726 255218 262210 255454
rect 262446 255218 292930 255454
rect 293166 255218 323650 255454
rect 323886 255218 354370 255454
rect 354606 255218 385090 255454
rect 385326 255218 415810 255454
rect 416046 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 586890 255454
rect -2966 255134 586890 255218
rect -2966 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 73826 255134
rect 74062 254898 74146 255134
rect 74382 254898 109826 255134
rect 110062 254898 110146 255134
rect 110382 254898 145826 255134
rect 146062 254898 146146 255134
rect 146382 254898 170050 255134
rect 170286 254898 200770 255134
rect 201006 254898 231490 255134
rect 231726 254898 262210 255134
rect 262446 254898 292930 255134
rect 293166 254898 323650 255134
rect 323886 254898 354370 255134
rect 354606 254898 385090 255134
rect 385326 254898 415810 255134
rect 416046 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 586890 255134
rect -2966 254866 586890 254898
rect -8726 248614 592650 248646
rect -8726 248378 -8694 248614
rect -8458 248378 -8374 248614
rect -8138 248378 30986 248614
rect 31222 248378 31306 248614
rect 31542 248378 66986 248614
rect 67222 248378 67306 248614
rect 67542 248378 102986 248614
rect 103222 248378 103306 248614
rect 103542 248378 138986 248614
rect 139222 248378 139306 248614
rect 139542 248378 426986 248614
rect 427222 248378 427306 248614
rect 427542 248378 462986 248614
rect 463222 248378 463306 248614
rect 463542 248378 498986 248614
rect 499222 248378 499306 248614
rect 499542 248378 534986 248614
rect 535222 248378 535306 248614
rect 535542 248378 570986 248614
rect 571222 248378 571306 248614
rect 571542 248378 592062 248614
rect 592298 248378 592382 248614
rect 592618 248378 592650 248614
rect -8726 248294 592650 248378
rect -8726 248058 -8694 248294
rect -8458 248058 -8374 248294
rect -8138 248058 30986 248294
rect 31222 248058 31306 248294
rect 31542 248058 66986 248294
rect 67222 248058 67306 248294
rect 67542 248058 102986 248294
rect 103222 248058 103306 248294
rect 103542 248058 138986 248294
rect 139222 248058 139306 248294
rect 139542 248058 426986 248294
rect 427222 248058 427306 248294
rect 427542 248058 462986 248294
rect 463222 248058 463306 248294
rect 463542 248058 498986 248294
rect 499222 248058 499306 248294
rect 499542 248058 534986 248294
rect 535222 248058 535306 248294
rect 535542 248058 570986 248294
rect 571222 248058 571306 248294
rect 571542 248058 592062 248294
rect 592298 248058 592382 248294
rect 592618 248058 592650 248294
rect -8726 248026 592650 248058
rect -6806 244894 590730 244926
rect -6806 244658 -6774 244894
rect -6538 244658 -6454 244894
rect -6218 244658 27266 244894
rect 27502 244658 27586 244894
rect 27822 244658 63266 244894
rect 63502 244658 63586 244894
rect 63822 244658 99266 244894
rect 99502 244658 99586 244894
rect 99822 244658 135266 244894
rect 135502 244658 135586 244894
rect 135822 244658 423266 244894
rect 423502 244658 423586 244894
rect 423822 244658 459266 244894
rect 459502 244658 459586 244894
rect 459822 244658 495266 244894
rect 495502 244658 495586 244894
rect 495822 244658 531266 244894
rect 531502 244658 531586 244894
rect 531822 244658 567266 244894
rect 567502 244658 567586 244894
rect 567822 244658 590142 244894
rect 590378 244658 590462 244894
rect 590698 244658 590730 244894
rect -6806 244574 590730 244658
rect -6806 244338 -6774 244574
rect -6538 244338 -6454 244574
rect -6218 244338 27266 244574
rect 27502 244338 27586 244574
rect 27822 244338 63266 244574
rect 63502 244338 63586 244574
rect 63822 244338 99266 244574
rect 99502 244338 99586 244574
rect 99822 244338 135266 244574
rect 135502 244338 135586 244574
rect 135822 244338 423266 244574
rect 423502 244338 423586 244574
rect 423822 244338 459266 244574
rect 459502 244338 459586 244574
rect 459822 244338 495266 244574
rect 495502 244338 495586 244574
rect 495822 244338 531266 244574
rect 531502 244338 531586 244574
rect 531822 244338 567266 244574
rect 567502 244338 567586 244574
rect 567822 244338 590142 244574
rect 590378 244338 590462 244574
rect 590698 244338 590730 244574
rect -6806 244306 590730 244338
rect -4886 241174 588810 241206
rect -4886 240938 -4854 241174
rect -4618 240938 -4534 241174
rect -4298 240938 23546 241174
rect 23782 240938 23866 241174
rect 24102 240938 59546 241174
rect 59782 240938 59866 241174
rect 60102 240938 95546 241174
rect 95782 240938 95866 241174
rect 96102 240938 131546 241174
rect 131782 240938 131866 241174
rect 132102 240938 455546 241174
rect 455782 240938 455866 241174
rect 456102 240938 491546 241174
rect 491782 240938 491866 241174
rect 492102 240938 527546 241174
rect 527782 240938 527866 241174
rect 528102 240938 563546 241174
rect 563782 240938 563866 241174
rect 564102 240938 588222 241174
rect 588458 240938 588542 241174
rect 588778 240938 588810 241174
rect -4886 240854 588810 240938
rect -4886 240618 -4854 240854
rect -4618 240618 -4534 240854
rect -4298 240618 23546 240854
rect 23782 240618 23866 240854
rect 24102 240618 59546 240854
rect 59782 240618 59866 240854
rect 60102 240618 95546 240854
rect 95782 240618 95866 240854
rect 96102 240618 131546 240854
rect 131782 240618 131866 240854
rect 132102 240618 455546 240854
rect 455782 240618 455866 240854
rect 456102 240618 491546 240854
rect 491782 240618 491866 240854
rect 492102 240618 527546 240854
rect 527782 240618 527866 240854
rect 528102 240618 563546 240854
rect 563782 240618 563866 240854
rect 564102 240618 588222 240854
rect 588458 240618 588542 240854
rect 588778 240618 588810 240854
rect -4886 240586 588810 240618
rect -2966 237454 586890 237486
rect -2966 237218 -2934 237454
rect -2698 237218 -2614 237454
rect -2378 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 55826 237454
rect 56062 237218 56146 237454
rect 56382 237218 91826 237454
rect 92062 237218 92146 237454
rect 92382 237218 127826 237454
rect 128062 237218 128146 237454
rect 128382 237218 185410 237454
rect 185646 237218 216130 237454
rect 216366 237218 246850 237454
rect 247086 237218 277570 237454
rect 277806 237218 308290 237454
rect 308526 237218 339010 237454
rect 339246 237218 369730 237454
rect 369966 237218 400450 237454
rect 400686 237218 451826 237454
rect 452062 237218 452146 237454
rect 452382 237218 487826 237454
rect 488062 237218 488146 237454
rect 488382 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 586302 237454
rect 586538 237218 586622 237454
rect 586858 237218 586890 237454
rect -2966 237134 586890 237218
rect -2966 236898 -2934 237134
rect -2698 236898 -2614 237134
rect -2378 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 55826 237134
rect 56062 236898 56146 237134
rect 56382 236898 91826 237134
rect 92062 236898 92146 237134
rect 92382 236898 127826 237134
rect 128062 236898 128146 237134
rect 128382 236898 185410 237134
rect 185646 236898 216130 237134
rect 216366 236898 246850 237134
rect 247086 236898 277570 237134
rect 277806 236898 308290 237134
rect 308526 236898 339010 237134
rect 339246 236898 369730 237134
rect 369966 236898 400450 237134
rect 400686 236898 451826 237134
rect 452062 236898 452146 237134
rect 452382 236898 487826 237134
rect 488062 236898 488146 237134
rect 488382 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 586302 237134
rect 586538 236898 586622 237134
rect 586858 236898 586890 237134
rect -2966 236866 586890 236898
rect -8726 230614 592650 230646
rect -8726 230378 -7734 230614
rect -7498 230378 -7414 230614
rect -7178 230378 12986 230614
rect 13222 230378 13306 230614
rect 13542 230378 48986 230614
rect 49222 230378 49306 230614
rect 49542 230378 84986 230614
rect 85222 230378 85306 230614
rect 85542 230378 120986 230614
rect 121222 230378 121306 230614
rect 121542 230378 156986 230614
rect 157222 230378 157306 230614
rect 157542 230378 444986 230614
rect 445222 230378 445306 230614
rect 445542 230378 480986 230614
rect 481222 230378 481306 230614
rect 481542 230378 516986 230614
rect 517222 230378 517306 230614
rect 517542 230378 552986 230614
rect 553222 230378 553306 230614
rect 553542 230378 591102 230614
rect 591338 230378 591422 230614
rect 591658 230378 592650 230614
rect -8726 230294 592650 230378
rect -8726 230058 -7734 230294
rect -7498 230058 -7414 230294
rect -7178 230058 12986 230294
rect 13222 230058 13306 230294
rect 13542 230058 48986 230294
rect 49222 230058 49306 230294
rect 49542 230058 84986 230294
rect 85222 230058 85306 230294
rect 85542 230058 120986 230294
rect 121222 230058 121306 230294
rect 121542 230058 156986 230294
rect 157222 230058 157306 230294
rect 157542 230058 444986 230294
rect 445222 230058 445306 230294
rect 445542 230058 480986 230294
rect 481222 230058 481306 230294
rect 481542 230058 516986 230294
rect 517222 230058 517306 230294
rect 517542 230058 552986 230294
rect 553222 230058 553306 230294
rect 553542 230058 591102 230294
rect 591338 230058 591422 230294
rect 591658 230058 592650 230294
rect -8726 230026 592650 230058
rect -6806 226894 590730 226926
rect -6806 226658 -5814 226894
rect -5578 226658 -5494 226894
rect -5258 226658 9266 226894
rect 9502 226658 9586 226894
rect 9822 226658 45266 226894
rect 45502 226658 45586 226894
rect 45822 226658 81266 226894
rect 81502 226658 81586 226894
rect 81822 226658 117266 226894
rect 117502 226658 117586 226894
rect 117822 226658 153266 226894
rect 153502 226658 153586 226894
rect 153822 226658 441266 226894
rect 441502 226658 441586 226894
rect 441822 226658 477266 226894
rect 477502 226658 477586 226894
rect 477822 226658 513266 226894
rect 513502 226658 513586 226894
rect 513822 226658 549266 226894
rect 549502 226658 549586 226894
rect 549822 226658 589182 226894
rect 589418 226658 589502 226894
rect 589738 226658 590730 226894
rect -6806 226574 590730 226658
rect -6806 226338 -5814 226574
rect -5578 226338 -5494 226574
rect -5258 226338 9266 226574
rect 9502 226338 9586 226574
rect 9822 226338 45266 226574
rect 45502 226338 45586 226574
rect 45822 226338 81266 226574
rect 81502 226338 81586 226574
rect 81822 226338 117266 226574
rect 117502 226338 117586 226574
rect 117822 226338 153266 226574
rect 153502 226338 153586 226574
rect 153822 226338 441266 226574
rect 441502 226338 441586 226574
rect 441822 226338 477266 226574
rect 477502 226338 477586 226574
rect 477822 226338 513266 226574
rect 513502 226338 513586 226574
rect 513822 226338 549266 226574
rect 549502 226338 549586 226574
rect 549822 226338 589182 226574
rect 589418 226338 589502 226574
rect 589738 226338 590730 226574
rect -6806 226306 590730 226338
rect -4886 223174 588810 223206
rect -4886 222938 -3894 223174
rect -3658 222938 -3574 223174
rect -3338 222938 5546 223174
rect 5782 222938 5866 223174
rect 6102 222938 41546 223174
rect 41782 222938 41866 223174
rect 42102 222938 77546 223174
rect 77782 222938 77866 223174
rect 78102 222938 113546 223174
rect 113782 222938 113866 223174
rect 114102 222938 149546 223174
rect 149782 222938 149866 223174
rect 150102 222938 437546 223174
rect 437782 222938 437866 223174
rect 438102 222938 473546 223174
rect 473782 222938 473866 223174
rect 474102 222938 509546 223174
rect 509782 222938 509866 223174
rect 510102 222938 545546 223174
rect 545782 222938 545866 223174
rect 546102 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 587262 223174
rect 587498 222938 587582 223174
rect 587818 222938 588810 223174
rect -4886 222854 588810 222938
rect -4886 222618 -3894 222854
rect -3658 222618 -3574 222854
rect -3338 222618 5546 222854
rect 5782 222618 5866 222854
rect 6102 222618 41546 222854
rect 41782 222618 41866 222854
rect 42102 222618 77546 222854
rect 77782 222618 77866 222854
rect 78102 222618 113546 222854
rect 113782 222618 113866 222854
rect 114102 222618 149546 222854
rect 149782 222618 149866 222854
rect 150102 222618 437546 222854
rect 437782 222618 437866 222854
rect 438102 222618 473546 222854
rect 473782 222618 473866 222854
rect 474102 222618 509546 222854
rect 509782 222618 509866 222854
rect 510102 222618 545546 222854
rect 545782 222618 545866 222854
rect 546102 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 587262 222854
rect 587498 222618 587582 222854
rect 587818 222618 588810 222854
rect -4886 222586 588810 222618
rect -2966 219454 586890 219486
rect -2966 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 73826 219454
rect 74062 219218 74146 219454
rect 74382 219218 109826 219454
rect 110062 219218 110146 219454
rect 110382 219218 145826 219454
rect 146062 219218 146146 219454
rect 146382 219218 170050 219454
rect 170286 219218 200770 219454
rect 201006 219218 231490 219454
rect 231726 219218 262210 219454
rect 262446 219218 292930 219454
rect 293166 219218 323650 219454
rect 323886 219218 354370 219454
rect 354606 219218 385090 219454
rect 385326 219218 415810 219454
rect 416046 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 586890 219454
rect -2966 219134 586890 219218
rect -2966 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 73826 219134
rect 74062 218898 74146 219134
rect 74382 218898 109826 219134
rect 110062 218898 110146 219134
rect 110382 218898 145826 219134
rect 146062 218898 146146 219134
rect 146382 218898 170050 219134
rect 170286 218898 200770 219134
rect 201006 218898 231490 219134
rect 231726 218898 262210 219134
rect 262446 218898 292930 219134
rect 293166 218898 323650 219134
rect 323886 218898 354370 219134
rect 354606 218898 385090 219134
rect 385326 218898 415810 219134
rect 416046 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 586890 219134
rect -2966 218866 586890 218898
rect -8726 212614 592650 212646
rect -8726 212378 -8694 212614
rect -8458 212378 -8374 212614
rect -8138 212378 30986 212614
rect 31222 212378 31306 212614
rect 31542 212378 66986 212614
rect 67222 212378 67306 212614
rect 67542 212378 102986 212614
rect 103222 212378 103306 212614
rect 103542 212378 138986 212614
rect 139222 212378 139306 212614
rect 139542 212378 426986 212614
rect 427222 212378 427306 212614
rect 427542 212378 462986 212614
rect 463222 212378 463306 212614
rect 463542 212378 498986 212614
rect 499222 212378 499306 212614
rect 499542 212378 534986 212614
rect 535222 212378 535306 212614
rect 535542 212378 570986 212614
rect 571222 212378 571306 212614
rect 571542 212378 592062 212614
rect 592298 212378 592382 212614
rect 592618 212378 592650 212614
rect -8726 212294 592650 212378
rect -8726 212058 -8694 212294
rect -8458 212058 -8374 212294
rect -8138 212058 30986 212294
rect 31222 212058 31306 212294
rect 31542 212058 66986 212294
rect 67222 212058 67306 212294
rect 67542 212058 102986 212294
rect 103222 212058 103306 212294
rect 103542 212058 138986 212294
rect 139222 212058 139306 212294
rect 139542 212058 426986 212294
rect 427222 212058 427306 212294
rect 427542 212058 462986 212294
rect 463222 212058 463306 212294
rect 463542 212058 498986 212294
rect 499222 212058 499306 212294
rect 499542 212058 534986 212294
rect 535222 212058 535306 212294
rect 535542 212058 570986 212294
rect 571222 212058 571306 212294
rect 571542 212058 592062 212294
rect 592298 212058 592382 212294
rect 592618 212058 592650 212294
rect -8726 212026 592650 212058
rect -6806 208894 590730 208926
rect -6806 208658 -6774 208894
rect -6538 208658 -6454 208894
rect -6218 208658 27266 208894
rect 27502 208658 27586 208894
rect 27822 208658 63266 208894
rect 63502 208658 63586 208894
rect 63822 208658 99266 208894
rect 99502 208658 99586 208894
rect 99822 208658 135266 208894
rect 135502 208658 135586 208894
rect 135822 208658 423266 208894
rect 423502 208658 423586 208894
rect 423822 208658 459266 208894
rect 459502 208658 459586 208894
rect 459822 208658 495266 208894
rect 495502 208658 495586 208894
rect 495822 208658 531266 208894
rect 531502 208658 531586 208894
rect 531822 208658 567266 208894
rect 567502 208658 567586 208894
rect 567822 208658 590142 208894
rect 590378 208658 590462 208894
rect 590698 208658 590730 208894
rect -6806 208574 590730 208658
rect -6806 208338 -6774 208574
rect -6538 208338 -6454 208574
rect -6218 208338 27266 208574
rect 27502 208338 27586 208574
rect 27822 208338 63266 208574
rect 63502 208338 63586 208574
rect 63822 208338 99266 208574
rect 99502 208338 99586 208574
rect 99822 208338 135266 208574
rect 135502 208338 135586 208574
rect 135822 208338 423266 208574
rect 423502 208338 423586 208574
rect 423822 208338 459266 208574
rect 459502 208338 459586 208574
rect 459822 208338 495266 208574
rect 495502 208338 495586 208574
rect 495822 208338 531266 208574
rect 531502 208338 531586 208574
rect 531822 208338 567266 208574
rect 567502 208338 567586 208574
rect 567822 208338 590142 208574
rect 590378 208338 590462 208574
rect 590698 208338 590730 208574
rect -6806 208306 590730 208338
rect -4886 205174 588810 205206
rect -4886 204938 -4854 205174
rect -4618 204938 -4534 205174
rect -4298 204938 23546 205174
rect 23782 204938 23866 205174
rect 24102 204938 59546 205174
rect 59782 204938 59866 205174
rect 60102 204938 95546 205174
rect 95782 204938 95866 205174
rect 96102 204938 131546 205174
rect 131782 204938 131866 205174
rect 132102 204938 455546 205174
rect 455782 204938 455866 205174
rect 456102 204938 491546 205174
rect 491782 204938 491866 205174
rect 492102 204938 527546 205174
rect 527782 204938 527866 205174
rect 528102 204938 563546 205174
rect 563782 204938 563866 205174
rect 564102 204938 588222 205174
rect 588458 204938 588542 205174
rect 588778 204938 588810 205174
rect -4886 204854 588810 204938
rect -4886 204618 -4854 204854
rect -4618 204618 -4534 204854
rect -4298 204618 23546 204854
rect 23782 204618 23866 204854
rect 24102 204618 59546 204854
rect 59782 204618 59866 204854
rect 60102 204618 95546 204854
rect 95782 204618 95866 204854
rect 96102 204618 131546 204854
rect 131782 204618 131866 204854
rect 132102 204618 455546 204854
rect 455782 204618 455866 204854
rect 456102 204618 491546 204854
rect 491782 204618 491866 204854
rect 492102 204618 527546 204854
rect 527782 204618 527866 204854
rect 528102 204618 563546 204854
rect 563782 204618 563866 204854
rect 564102 204618 588222 204854
rect 588458 204618 588542 204854
rect 588778 204618 588810 204854
rect -4886 204586 588810 204618
rect -2966 201454 586890 201486
rect -2966 201218 -2934 201454
rect -2698 201218 -2614 201454
rect -2378 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 91826 201454
rect 92062 201218 92146 201454
rect 92382 201218 127826 201454
rect 128062 201218 128146 201454
rect 128382 201218 451826 201454
rect 452062 201218 452146 201454
rect 452382 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 586302 201454
rect 586538 201218 586622 201454
rect 586858 201218 586890 201454
rect -2966 201134 586890 201218
rect -2966 200898 -2934 201134
rect -2698 200898 -2614 201134
rect -2378 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 91826 201134
rect 92062 200898 92146 201134
rect 92382 200898 127826 201134
rect 128062 200898 128146 201134
rect 128382 200898 451826 201134
rect 452062 200898 452146 201134
rect 452382 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 586302 201134
rect 586538 200898 586622 201134
rect 586858 200898 586890 201134
rect -2966 200866 586890 200898
rect -8726 194614 592650 194646
rect -8726 194378 -7734 194614
rect -7498 194378 -7414 194614
rect -7178 194378 12986 194614
rect 13222 194378 13306 194614
rect 13542 194378 48986 194614
rect 49222 194378 49306 194614
rect 49542 194378 84986 194614
rect 85222 194378 85306 194614
rect 85542 194378 120986 194614
rect 121222 194378 121306 194614
rect 121542 194378 156986 194614
rect 157222 194378 157306 194614
rect 157542 194378 192986 194614
rect 193222 194378 193306 194614
rect 193542 194378 228986 194614
rect 229222 194378 229306 194614
rect 229542 194378 264986 194614
rect 265222 194378 265306 194614
rect 265542 194378 300986 194614
rect 301222 194378 301306 194614
rect 301542 194378 336986 194614
rect 337222 194378 337306 194614
rect 337542 194378 372986 194614
rect 373222 194378 373306 194614
rect 373542 194378 408986 194614
rect 409222 194378 409306 194614
rect 409542 194378 444986 194614
rect 445222 194378 445306 194614
rect 445542 194378 480986 194614
rect 481222 194378 481306 194614
rect 481542 194378 516986 194614
rect 517222 194378 517306 194614
rect 517542 194378 552986 194614
rect 553222 194378 553306 194614
rect 553542 194378 591102 194614
rect 591338 194378 591422 194614
rect 591658 194378 592650 194614
rect -8726 194294 592650 194378
rect -8726 194058 -7734 194294
rect -7498 194058 -7414 194294
rect -7178 194058 12986 194294
rect 13222 194058 13306 194294
rect 13542 194058 48986 194294
rect 49222 194058 49306 194294
rect 49542 194058 84986 194294
rect 85222 194058 85306 194294
rect 85542 194058 120986 194294
rect 121222 194058 121306 194294
rect 121542 194058 156986 194294
rect 157222 194058 157306 194294
rect 157542 194058 192986 194294
rect 193222 194058 193306 194294
rect 193542 194058 228986 194294
rect 229222 194058 229306 194294
rect 229542 194058 264986 194294
rect 265222 194058 265306 194294
rect 265542 194058 300986 194294
rect 301222 194058 301306 194294
rect 301542 194058 336986 194294
rect 337222 194058 337306 194294
rect 337542 194058 372986 194294
rect 373222 194058 373306 194294
rect 373542 194058 408986 194294
rect 409222 194058 409306 194294
rect 409542 194058 444986 194294
rect 445222 194058 445306 194294
rect 445542 194058 480986 194294
rect 481222 194058 481306 194294
rect 481542 194058 516986 194294
rect 517222 194058 517306 194294
rect 517542 194058 552986 194294
rect 553222 194058 553306 194294
rect 553542 194058 591102 194294
rect 591338 194058 591422 194294
rect 591658 194058 592650 194294
rect -8726 194026 592650 194058
rect -6806 190894 590730 190926
rect -6806 190658 -5814 190894
rect -5578 190658 -5494 190894
rect -5258 190658 9266 190894
rect 9502 190658 9586 190894
rect 9822 190658 45266 190894
rect 45502 190658 45586 190894
rect 45822 190658 81266 190894
rect 81502 190658 81586 190894
rect 81822 190658 117266 190894
rect 117502 190658 117586 190894
rect 117822 190658 153266 190894
rect 153502 190658 153586 190894
rect 153822 190658 189266 190894
rect 189502 190658 189586 190894
rect 189822 190658 225266 190894
rect 225502 190658 225586 190894
rect 225822 190658 261266 190894
rect 261502 190658 261586 190894
rect 261822 190658 297266 190894
rect 297502 190658 297586 190894
rect 297822 190658 333266 190894
rect 333502 190658 333586 190894
rect 333822 190658 369266 190894
rect 369502 190658 369586 190894
rect 369822 190658 405266 190894
rect 405502 190658 405586 190894
rect 405822 190658 441266 190894
rect 441502 190658 441586 190894
rect 441822 190658 477266 190894
rect 477502 190658 477586 190894
rect 477822 190658 513266 190894
rect 513502 190658 513586 190894
rect 513822 190658 549266 190894
rect 549502 190658 549586 190894
rect 549822 190658 589182 190894
rect 589418 190658 589502 190894
rect 589738 190658 590730 190894
rect -6806 190574 590730 190658
rect -6806 190338 -5814 190574
rect -5578 190338 -5494 190574
rect -5258 190338 9266 190574
rect 9502 190338 9586 190574
rect 9822 190338 45266 190574
rect 45502 190338 45586 190574
rect 45822 190338 81266 190574
rect 81502 190338 81586 190574
rect 81822 190338 117266 190574
rect 117502 190338 117586 190574
rect 117822 190338 153266 190574
rect 153502 190338 153586 190574
rect 153822 190338 189266 190574
rect 189502 190338 189586 190574
rect 189822 190338 225266 190574
rect 225502 190338 225586 190574
rect 225822 190338 261266 190574
rect 261502 190338 261586 190574
rect 261822 190338 297266 190574
rect 297502 190338 297586 190574
rect 297822 190338 333266 190574
rect 333502 190338 333586 190574
rect 333822 190338 369266 190574
rect 369502 190338 369586 190574
rect 369822 190338 405266 190574
rect 405502 190338 405586 190574
rect 405822 190338 441266 190574
rect 441502 190338 441586 190574
rect 441822 190338 477266 190574
rect 477502 190338 477586 190574
rect 477822 190338 513266 190574
rect 513502 190338 513586 190574
rect 513822 190338 549266 190574
rect 549502 190338 549586 190574
rect 549822 190338 589182 190574
rect 589418 190338 589502 190574
rect 589738 190338 590730 190574
rect -6806 190306 590730 190338
rect -4886 187174 588810 187206
rect -4886 186938 -3894 187174
rect -3658 186938 -3574 187174
rect -3338 186938 5546 187174
rect 5782 186938 5866 187174
rect 6102 186938 41546 187174
rect 41782 186938 41866 187174
rect 42102 186938 77546 187174
rect 77782 186938 77866 187174
rect 78102 186938 113546 187174
rect 113782 186938 113866 187174
rect 114102 186938 149546 187174
rect 149782 186938 149866 187174
rect 150102 186938 185546 187174
rect 185782 186938 185866 187174
rect 186102 186938 221546 187174
rect 221782 186938 221866 187174
rect 222102 186938 257546 187174
rect 257782 186938 257866 187174
rect 258102 186938 293546 187174
rect 293782 186938 293866 187174
rect 294102 186938 329546 187174
rect 329782 186938 329866 187174
rect 330102 186938 365546 187174
rect 365782 186938 365866 187174
rect 366102 186938 401546 187174
rect 401782 186938 401866 187174
rect 402102 186938 437546 187174
rect 437782 186938 437866 187174
rect 438102 186938 473546 187174
rect 473782 186938 473866 187174
rect 474102 186938 509546 187174
rect 509782 186938 509866 187174
rect 510102 186938 545546 187174
rect 545782 186938 545866 187174
rect 546102 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 587262 187174
rect 587498 186938 587582 187174
rect 587818 186938 588810 187174
rect -4886 186854 588810 186938
rect -4886 186618 -3894 186854
rect -3658 186618 -3574 186854
rect -3338 186618 5546 186854
rect 5782 186618 5866 186854
rect 6102 186618 41546 186854
rect 41782 186618 41866 186854
rect 42102 186618 77546 186854
rect 77782 186618 77866 186854
rect 78102 186618 113546 186854
rect 113782 186618 113866 186854
rect 114102 186618 149546 186854
rect 149782 186618 149866 186854
rect 150102 186618 185546 186854
rect 185782 186618 185866 186854
rect 186102 186618 221546 186854
rect 221782 186618 221866 186854
rect 222102 186618 257546 186854
rect 257782 186618 257866 186854
rect 258102 186618 293546 186854
rect 293782 186618 293866 186854
rect 294102 186618 329546 186854
rect 329782 186618 329866 186854
rect 330102 186618 365546 186854
rect 365782 186618 365866 186854
rect 366102 186618 401546 186854
rect 401782 186618 401866 186854
rect 402102 186618 437546 186854
rect 437782 186618 437866 186854
rect 438102 186618 473546 186854
rect 473782 186618 473866 186854
rect 474102 186618 509546 186854
rect 509782 186618 509866 186854
rect 510102 186618 545546 186854
rect 545782 186618 545866 186854
rect 546102 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 587262 186854
rect 587498 186618 587582 186854
rect 587818 186618 588810 186854
rect -4886 186586 588810 186618
rect -2966 183454 586890 183486
rect -2966 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 73826 183454
rect 74062 183218 74146 183454
rect 74382 183218 109826 183454
rect 110062 183218 110146 183454
rect 110382 183218 145826 183454
rect 146062 183218 146146 183454
rect 146382 183218 181826 183454
rect 182062 183218 182146 183454
rect 182382 183218 217826 183454
rect 218062 183218 218146 183454
rect 218382 183218 253826 183454
rect 254062 183218 254146 183454
rect 254382 183218 289826 183454
rect 290062 183218 290146 183454
rect 290382 183218 325826 183454
rect 326062 183218 326146 183454
rect 326382 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 586890 183454
rect -2966 183134 586890 183218
rect -2966 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 73826 183134
rect 74062 182898 74146 183134
rect 74382 182898 109826 183134
rect 110062 182898 110146 183134
rect 110382 182898 145826 183134
rect 146062 182898 146146 183134
rect 146382 182898 181826 183134
rect 182062 182898 182146 183134
rect 182382 182898 217826 183134
rect 218062 182898 218146 183134
rect 218382 182898 253826 183134
rect 254062 182898 254146 183134
rect 254382 182898 289826 183134
rect 290062 182898 290146 183134
rect 290382 182898 325826 183134
rect 326062 182898 326146 183134
rect 326382 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 586890 183134
rect -2966 182866 586890 182898
rect -8726 176614 592650 176646
rect -8726 176378 -8694 176614
rect -8458 176378 -8374 176614
rect -8138 176378 30986 176614
rect 31222 176378 31306 176614
rect 31542 176378 66986 176614
rect 67222 176378 67306 176614
rect 67542 176378 102986 176614
rect 103222 176378 103306 176614
rect 103542 176378 138986 176614
rect 139222 176378 139306 176614
rect 139542 176378 174986 176614
rect 175222 176378 175306 176614
rect 175542 176378 210986 176614
rect 211222 176378 211306 176614
rect 211542 176378 246986 176614
rect 247222 176378 247306 176614
rect 247542 176378 282986 176614
rect 283222 176378 283306 176614
rect 283542 176378 318986 176614
rect 319222 176378 319306 176614
rect 319542 176378 354986 176614
rect 355222 176378 355306 176614
rect 355542 176378 390986 176614
rect 391222 176378 391306 176614
rect 391542 176378 426986 176614
rect 427222 176378 427306 176614
rect 427542 176378 462986 176614
rect 463222 176378 463306 176614
rect 463542 176378 498986 176614
rect 499222 176378 499306 176614
rect 499542 176378 534986 176614
rect 535222 176378 535306 176614
rect 535542 176378 570986 176614
rect 571222 176378 571306 176614
rect 571542 176378 592062 176614
rect 592298 176378 592382 176614
rect 592618 176378 592650 176614
rect -8726 176294 592650 176378
rect -8726 176058 -8694 176294
rect -8458 176058 -8374 176294
rect -8138 176058 30986 176294
rect 31222 176058 31306 176294
rect 31542 176058 66986 176294
rect 67222 176058 67306 176294
rect 67542 176058 102986 176294
rect 103222 176058 103306 176294
rect 103542 176058 138986 176294
rect 139222 176058 139306 176294
rect 139542 176058 174986 176294
rect 175222 176058 175306 176294
rect 175542 176058 210986 176294
rect 211222 176058 211306 176294
rect 211542 176058 246986 176294
rect 247222 176058 247306 176294
rect 247542 176058 282986 176294
rect 283222 176058 283306 176294
rect 283542 176058 318986 176294
rect 319222 176058 319306 176294
rect 319542 176058 354986 176294
rect 355222 176058 355306 176294
rect 355542 176058 390986 176294
rect 391222 176058 391306 176294
rect 391542 176058 426986 176294
rect 427222 176058 427306 176294
rect 427542 176058 462986 176294
rect 463222 176058 463306 176294
rect 463542 176058 498986 176294
rect 499222 176058 499306 176294
rect 499542 176058 534986 176294
rect 535222 176058 535306 176294
rect 535542 176058 570986 176294
rect 571222 176058 571306 176294
rect 571542 176058 592062 176294
rect 592298 176058 592382 176294
rect 592618 176058 592650 176294
rect -8726 176026 592650 176058
rect -6806 172894 590730 172926
rect -6806 172658 -6774 172894
rect -6538 172658 -6454 172894
rect -6218 172658 27266 172894
rect 27502 172658 27586 172894
rect 27822 172658 63266 172894
rect 63502 172658 63586 172894
rect 63822 172658 99266 172894
rect 99502 172658 99586 172894
rect 99822 172658 135266 172894
rect 135502 172658 135586 172894
rect 135822 172658 171266 172894
rect 171502 172658 171586 172894
rect 171822 172658 207266 172894
rect 207502 172658 207586 172894
rect 207822 172658 243266 172894
rect 243502 172658 243586 172894
rect 243822 172658 279266 172894
rect 279502 172658 279586 172894
rect 279822 172658 315266 172894
rect 315502 172658 315586 172894
rect 315822 172658 351266 172894
rect 351502 172658 351586 172894
rect 351822 172658 387266 172894
rect 387502 172658 387586 172894
rect 387822 172658 423266 172894
rect 423502 172658 423586 172894
rect 423822 172658 459266 172894
rect 459502 172658 459586 172894
rect 459822 172658 495266 172894
rect 495502 172658 495586 172894
rect 495822 172658 531266 172894
rect 531502 172658 531586 172894
rect 531822 172658 567266 172894
rect 567502 172658 567586 172894
rect 567822 172658 590142 172894
rect 590378 172658 590462 172894
rect 590698 172658 590730 172894
rect -6806 172574 590730 172658
rect -6806 172338 -6774 172574
rect -6538 172338 -6454 172574
rect -6218 172338 27266 172574
rect 27502 172338 27586 172574
rect 27822 172338 63266 172574
rect 63502 172338 63586 172574
rect 63822 172338 99266 172574
rect 99502 172338 99586 172574
rect 99822 172338 135266 172574
rect 135502 172338 135586 172574
rect 135822 172338 171266 172574
rect 171502 172338 171586 172574
rect 171822 172338 207266 172574
rect 207502 172338 207586 172574
rect 207822 172338 243266 172574
rect 243502 172338 243586 172574
rect 243822 172338 279266 172574
rect 279502 172338 279586 172574
rect 279822 172338 315266 172574
rect 315502 172338 315586 172574
rect 315822 172338 351266 172574
rect 351502 172338 351586 172574
rect 351822 172338 387266 172574
rect 387502 172338 387586 172574
rect 387822 172338 423266 172574
rect 423502 172338 423586 172574
rect 423822 172338 459266 172574
rect 459502 172338 459586 172574
rect 459822 172338 495266 172574
rect 495502 172338 495586 172574
rect 495822 172338 531266 172574
rect 531502 172338 531586 172574
rect 531822 172338 567266 172574
rect 567502 172338 567586 172574
rect 567822 172338 590142 172574
rect 590378 172338 590462 172574
rect 590698 172338 590730 172574
rect -6806 172306 590730 172338
rect -4886 169174 588810 169206
rect -4886 168938 -4854 169174
rect -4618 168938 -4534 169174
rect -4298 168938 23546 169174
rect 23782 168938 23866 169174
rect 24102 168938 59546 169174
rect 59782 168938 59866 169174
rect 60102 168938 95546 169174
rect 95782 168938 95866 169174
rect 96102 168938 131546 169174
rect 131782 168938 131866 169174
rect 132102 168938 167546 169174
rect 167782 168938 167866 169174
rect 168102 168938 203546 169174
rect 203782 168938 203866 169174
rect 204102 168938 239546 169174
rect 239782 168938 239866 169174
rect 240102 168938 275546 169174
rect 275782 168938 275866 169174
rect 276102 168938 311546 169174
rect 311782 168938 311866 169174
rect 312102 168938 347546 169174
rect 347782 168938 347866 169174
rect 348102 168938 383546 169174
rect 383782 168938 383866 169174
rect 384102 168938 419546 169174
rect 419782 168938 419866 169174
rect 420102 168938 455546 169174
rect 455782 168938 455866 169174
rect 456102 168938 491546 169174
rect 491782 168938 491866 169174
rect 492102 168938 527546 169174
rect 527782 168938 527866 169174
rect 528102 168938 563546 169174
rect 563782 168938 563866 169174
rect 564102 168938 588222 169174
rect 588458 168938 588542 169174
rect 588778 168938 588810 169174
rect -4886 168854 588810 168938
rect -4886 168618 -4854 168854
rect -4618 168618 -4534 168854
rect -4298 168618 23546 168854
rect 23782 168618 23866 168854
rect 24102 168618 59546 168854
rect 59782 168618 59866 168854
rect 60102 168618 95546 168854
rect 95782 168618 95866 168854
rect 96102 168618 131546 168854
rect 131782 168618 131866 168854
rect 132102 168618 167546 168854
rect 167782 168618 167866 168854
rect 168102 168618 203546 168854
rect 203782 168618 203866 168854
rect 204102 168618 239546 168854
rect 239782 168618 239866 168854
rect 240102 168618 275546 168854
rect 275782 168618 275866 168854
rect 276102 168618 311546 168854
rect 311782 168618 311866 168854
rect 312102 168618 347546 168854
rect 347782 168618 347866 168854
rect 348102 168618 383546 168854
rect 383782 168618 383866 168854
rect 384102 168618 419546 168854
rect 419782 168618 419866 168854
rect 420102 168618 455546 168854
rect 455782 168618 455866 168854
rect 456102 168618 491546 168854
rect 491782 168618 491866 168854
rect 492102 168618 527546 168854
rect 527782 168618 527866 168854
rect 528102 168618 563546 168854
rect 563782 168618 563866 168854
rect 564102 168618 588222 168854
rect 588458 168618 588542 168854
rect 588778 168618 588810 168854
rect -4886 168586 588810 168618
rect -2966 165454 586890 165486
rect -2966 165218 -2934 165454
rect -2698 165218 -2614 165454
rect -2378 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 91826 165454
rect 92062 165218 92146 165454
rect 92382 165218 127826 165454
rect 128062 165218 128146 165454
rect 128382 165218 163826 165454
rect 164062 165218 164146 165454
rect 164382 165218 199826 165454
rect 200062 165218 200146 165454
rect 200382 165218 235826 165454
rect 236062 165218 236146 165454
rect 236382 165218 271826 165454
rect 272062 165218 272146 165454
rect 272382 165218 307826 165454
rect 308062 165218 308146 165454
rect 308382 165218 343826 165454
rect 344062 165218 344146 165454
rect 344382 165218 379826 165454
rect 380062 165218 380146 165454
rect 380382 165218 415826 165454
rect 416062 165218 416146 165454
rect 416382 165218 451826 165454
rect 452062 165218 452146 165454
rect 452382 165218 487826 165454
rect 488062 165218 488146 165454
rect 488382 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 586302 165454
rect 586538 165218 586622 165454
rect 586858 165218 586890 165454
rect -2966 165134 586890 165218
rect -2966 164898 -2934 165134
rect -2698 164898 -2614 165134
rect -2378 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 91826 165134
rect 92062 164898 92146 165134
rect 92382 164898 127826 165134
rect 128062 164898 128146 165134
rect 128382 164898 163826 165134
rect 164062 164898 164146 165134
rect 164382 164898 199826 165134
rect 200062 164898 200146 165134
rect 200382 164898 235826 165134
rect 236062 164898 236146 165134
rect 236382 164898 271826 165134
rect 272062 164898 272146 165134
rect 272382 164898 307826 165134
rect 308062 164898 308146 165134
rect 308382 164898 343826 165134
rect 344062 164898 344146 165134
rect 344382 164898 379826 165134
rect 380062 164898 380146 165134
rect 380382 164898 415826 165134
rect 416062 164898 416146 165134
rect 416382 164898 451826 165134
rect 452062 164898 452146 165134
rect 452382 164898 487826 165134
rect 488062 164898 488146 165134
rect 488382 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 586302 165134
rect 586538 164898 586622 165134
rect 586858 164898 586890 165134
rect -2966 164866 586890 164898
rect -8726 158614 592650 158646
rect -8726 158378 -7734 158614
rect -7498 158378 -7414 158614
rect -7178 158378 12986 158614
rect 13222 158378 13306 158614
rect 13542 158378 48986 158614
rect 49222 158378 49306 158614
rect 49542 158378 84986 158614
rect 85222 158378 85306 158614
rect 85542 158378 120986 158614
rect 121222 158378 121306 158614
rect 121542 158378 156986 158614
rect 157222 158378 157306 158614
rect 157542 158378 192986 158614
rect 193222 158378 193306 158614
rect 193542 158378 228986 158614
rect 229222 158378 229306 158614
rect 229542 158378 264986 158614
rect 265222 158378 265306 158614
rect 265542 158378 300986 158614
rect 301222 158378 301306 158614
rect 301542 158378 336986 158614
rect 337222 158378 337306 158614
rect 337542 158378 372986 158614
rect 373222 158378 373306 158614
rect 373542 158378 408986 158614
rect 409222 158378 409306 158614
rect 409542 158378 444986 158614
rect 445222 158378 445306 158614
rect 445542 158378 480986 158614
rect 481222 158378 481306 158614
rect 481542 158378 516986 158614
rect 517222 158378 517306 158614
rect 517542 158378 552986 158614
rect 553222 158378 553306 158614
rect 553542 158378 591102 158614
rect 591338 158378 591422 158614
rect 591658 158378 592650 158614
rect -8726 158294 592650 158378
rect -8726 158058 -7734 158294
rect -7498 158058 -7414 158294
rect -7178 158058 12986 158294
rect 13222 158058 13306 158294
rect 13542 158058 48986 158294
rect 49222 158058 49306 158294
rect 49542 158058 84986 158294
rect 85222 158058 85306 158294
rect 85542 158058 120986 158294
rect 121222 158058 121306 158294
rect 121542 158058 156986 158294
rect 157222 158058 157306 158294
rect 157542 158058 192986 158294
rect 193222 158058 193306 158294
rect 193542 158058 228986 158294
rect 229222 158058 229306 158294
rect 229542 158058 264986 158294
rect 265222 158058 265306 158294
rect 265542 158058 300986 158294
rect 301222 158058 301306 158294
rect 301542 158058 336986 158294
rect 337222 158058 337306 158294
rect 337542 158058 372986 158294
rect 373222 158058 373306 158294
rect 373542 158058 408986 158294
rect 409222 158058 409306 158294
rect 409542 158058 444986 158294
rect 445222 158058 445306 158294
rect 445542 158058 480986 158294
rect 481222 158058 481306 158294
rect 481542 158058 516986 158294
rect 517222 158058 517306 158294
rect 517542 158058 552986 158294
rect 553222 158058 553306 158294
rect 553542 158058 591102 158294
rect 591338 158058 591422 158294
rect 591658 158058 592650 158294
rect -8726 158026 592650 158058
rect -6806 154894 590730 154926
rect -6806 154658 -5814 154894
rect -5578 154658 -5494 154894
rect -5258 154658 9266 154894
rect 9502 154658 9586 154894
rect 9822 154658 45266 154894
rect 45502 154658 45586 154894
rect 45822 154658 81266 154894
rect 81502 154658 81586 154894
rect 81822 154658 117266 154894
rect 117502 154658 117586 154894
rect 117822 154658 153266 154894
rect 153502 154658 153586 154894
rect 153822 154658 189266 154894
rect 189502 154658 189586 154894
rect 189822 154658 225266 154894
rect 225502 154658 225586 154894
rect 225822 154658 261266 154894
rect 261502 154658 261586 154894
rect 261822 154658 297266 154894
rect 297502 154658 297586 154894
rect 297822 154658 333266 154894
rect 333502 154658 333586 154894
rect 333822 154658 369266 154894
rect 369502 154658 369586 154894
rect 369822 154658 405266 154894
rect 405502 154658 405586 154894
rect 405822 154658 441266 154894
rect 441502 154658 441586 154894
rect 441822 154658 477266 154894
rect 477502 154658 477586 154894
rect 477822 154658 513266 154894
rect 513502 154658 513586 154894
rect 513822 154658 549266 154894
rect 549502 154658 549586 154894
rect 549822 154658 589182 154894
rect 589418 154658 589502 154894
rect 589738 154658 590730 154894
rect -6806 154574 590730 154658
rect -6806 154338 -5814 154574
rect -5578 154338 -5494 154574
rect -5258 154338 9266 154574
rect 9502 154338 9586 154574
rect 9822 154338 45266 154574
rect 45502 154338 45586 154574
rect 45822 154338 81266 154574
rect 81502 154338 81586 154574
rect 81822 154338 117266 154574
rect 117502 154338 117586 154574
rect 117822 154338 153266 154574
rect 153502 154338 153586 154574
rect 153822 154338 189266 154574
rect 189502 154338 189586 154574
rect 189822 154338 225266 154574
rect 225502 154338 225586 154574
rect 225822 154338 261266 154574
rect 261502 154338 261586 154574
rect 261822 154338 297266 154574
rect 297502 154338 297586 154574
rect 297822 154338 333266 154574
rect 333502 154338 333586 154574
rect 333822 154338 369266 154574
rect 369502 154338 369586 154574
rect 369822 154338 405266 154574
rect 405502 154338 405586 154574
rect 405822 154338 441266 154574
rect 441502 154338 441586 154574
rect 441822 154338 477266 154574
rect 477502 154338 477586 154574
rect 477822 154338 513266 154574
rect 513502 154338 513586 154574
rect 513822 154338 549266 154574
rect 549502 154338 549586 154574
rect 549822 154338 589182 154574
rect 589418 154338 589502 154574
rect 589738 154338 590730 154574
rect -6806 154306 590730 154338
rect -4886 151174 588810 151206
rect -4886 150938 -3894 151174
rect -3658 150938 -3574 151174
rect -3338 150938 5546 151174
rect 5782 150938 5866 151174
rect 6102 150938 41546 151174
rect 41782 150938 41866 151174
rect 42102 150938 77546 151174
rect 77782 150938 77866 151174
rect 78102 150938 113546 151174
rect 113782 150938 113866 151174
rect 114102 150938 149546 151174
rect 149782 150938 149866 151174
rect 150102 150938 185546 151174
rect 185782 150938 185866 151174
rect 186102 150938 221546 151174
rect 221782 150938 221866 151174
rect 222102 150938 257546 151174
rect 257782 150938 257866 151174
rect 258102 150938 293546 151174
rect 293782 150938 293866 151174
rect 294102 150938 329546 151174
rect 329782 150938 329866 151174
rect 330102 150938 365546 151174
rect 365782 150938 365866 151174
rect 366102 150938 401546 151174
rect 401782 150938 401866 151174
rect 402102 150938 437546 151174
rect 437782 150938 437866 151174
rect 438102 150938 473546 151174
rect 473782 150938 473866 151174
rect 474102 150938 509546 151174
rect 509782 150938 509866 151174
rect 510102 150938 545546 151174
rect 545782 150938 545866 151174
rect 546102 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 587262 151174
rect 587498 150938 587582 151174
rect 587818 150938 588810 151174
rect -4886 150854 588810 150938
rect -4886 150618 -3894 150854
rect -3658 150618 -3574 150854
rect -3338 150618 5546 150854
rect 5782 150618 5866 150854
rect 6102 150618 41546 150854
rect 41782 150618 41866 150854
rect 42102 150618 77546 150854
rect 77782 150618 77866 150854
rect 78102 150618 113546 150854
rect 113782 150618 113866 150854
rect 114102 150618 149546 150854
rect 149782 150618 149866 150854
rect 150102 150618 185546 150854
rect 185782 150618 185866 150854
rect 186102 150618 221546 150854
rect 221782 150618 221866 150854
rect 222102 150618 257546 150854
rect 257782 150618 257866 150854
rect 258102 150618 293546 150854
rect 293782 150618 293866 150854
rect 294102 150618 329546 150854
rect 329782 150618 329866 150854
rect 330102 150618 365546 150854
rect 365782 150618 365866 150854
rect 366102 150618 401546 150854
rect 401782 150618 401866 150854
rect 402102 150618 437546 150854
rect 437782 150618 437866 150854
rect 438102 150618 473546 150854
rect 473782 150618 473866 150854
rect 474102 150618 509546 150854
rect 509782 150618 509866 150854
rect 510102 150618 545546 150854
rect 545782 150618 545866 150854
rect 546102 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 587262 150854
rect 587498 150618 587582 150854
rect 587818 150618 588810 150854
rect -4886 150586 588810 150618
rect -2966 147454 586890 147486
rect -2966 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 73826 147454
rect 74062 147218 74146 147454
rect 74382 147218 109826 147454
rect 110062 147218 110146 147454
rect 110382 147218 145826 147454
rect 146062 147218 146146 147454
rect 146382 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 217826 147454
rect 218062 147218 218146 147454
rect 218382 147218 253826 147454
rect 254062 147218 254146 147454
rect 254382 147218 289826 147454
rect 290062 147218 290146 147454
rect 290382 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 586890 147454
rect -2966 147134 586890 147218
rect -2966 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 73826 147134
rect 74062 146898 74146 147134
rect 74382 146898 109826 147134
rect 110062 146898 110146 147134
rect 110382 146898 145826 147134
rect 146062 146898 146146 147134
rect 146382 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 217826 147134
rect 218062 146898 218146 147134
rect 218382 146898 253826 147134
rect 254062 146898 254146 147134
rect 254382 146898 289826 147134
rect 290062 146898 290146 147134
rect 290382 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 586890 147134
rect -2966 146866 586890 146898
rect -8726 140614 592650 140646
rect -8726 140378 -8694 140614
rect -8458 140378 -8374 140614
rect -8138 140378 30986 140614
rect 31222 140378 31306 140614
rect 31542 140378 66986 140614
rect 67222 140378 67306 140614
rect 67542 140378 102986 140614
rect 103222 140378 103306 140614
rect 103542 140378 138986 140614
rect 139222 140378 139306 140614
rect 139542 140378 174986 140614
rect 175222 140378 175306 140614
rect 175542 140378 210986 140614
rect 211222 140378 211306 140614
rect 211542 140378 246986 140614
rect 247222 140378 247306 140614
rect 247542 140378 282986 140614
rect 283222 140378 283306 140614
rect 283542 140378 318986 140614
rect 319222 140378 319306 140614
rect 319542 140378 354986 140614
rect 355222 140378 355306 140614
rect 355542 140378 390986 140614
rect 391222 140378 391306 140614
rect 391542 140378 426986 140614
rect 427222 140378 427306 140614
rect 427542 140378 462986 140614
rect 463222 140378 463306 140614
rect 463542 140378 498986 140614
rect 499222 140378 499306 140614
rect 499542 140378 534986 140614
rect 535222 140378 535306 140614
rect 535542 140378 570986 140614
rect 571222 140378 571306 140614
rect 571542 140378 592062 140614
rect 592298 140378 592382 140614
rect 592618 140378 592650 140614
rect -8726 140294 592650 140378
rect -8726 140058 -8694 140294
rect -8458 140058 -8374 140294
rect -8138 140058 30986 140294
rect 31222 140058 31306 140294
rect 31542 140058 66986 140294
rect 67222 140058 67306 140294
rect 67542 140058 102986 140294
rect 103222 140058 103306 140294
rect 103542 140058 138986 140294
rect 139222 140058 139306 140294
rect 139542 140058 174986 140294
rect 175222 140058 175306 140294
rect 175542 140058 210986 140294
rect 211222 140058 211306 140294
rect 211542 140058 246986 140294
rect 247222 140058 247306 140294
rect 247542 140058 282986 140294
rect 283222 140058 283306 140294
rect 283542 140058 318986 140294
rect 319222 140058 319306 140294
rect 319542 140058 354986 140294
rect 355222 140058 355306 140294
rect 355542 140058 390986 140294
rect 391222 140058 391306 140294
rect 391542 140058 426986 140294
rect 427222 140058 427306 140294
rect 427542 140058 462986 140294
rect 463222 140058 463306 140294
rect 463542 140058 498986 140294
rect 499222 140058 499306 140294
rect 499542 140058 534986 140294
rect 535222 140058 535306 140294
rect 535542 140058 570986 140294
rect 571222 140058 571306 140294
rect 571542 140058 592062 140294
rect 592298 140058 592382 140294
rect 592618 140058 592650 140294
rect -8726 140026 592650 140058
rect -6806 136894 590730 136926
rect -6806 136658 -6774 136894
rect -6538 136658 -6454 136894
rect -6218 136658 27266 136894
rect 27502 136658 27586 136894
rect 27822 136658 63266 136894
rect 63502 136658 63586 136894
rect 63822 136658 99266 136894
rect 99502 136658 99586 136894
rect 99822 136658 135266 136894
rect 135502 136658 135586 136894
rect 135822 136658 171266 136894
rect 171502 136658 171586 136894
rect 171822 136658 207266 136894
rect 207502 136658 207586 136894
rect 207822 136658 243266 136894
rect 243502 136658 243586 136894
rect 243822 136658 279266 136894
rect 279502 136658 279586 136894
rect 279822 136658 315266 136894
rect 315502 136658 315586 136894
rect 315822 136658 351266 136894
rect 351502 136658 351586 136894
rect 351822 136658 387266 136894
rect 387502 136658 387586 136894
rect 387822 136658 423266 136894
rect 423502 136658 423586 136894
rect 423822 136658 459266 136894
rect 459502 136658 459586 136894
rect 459822 136658 495266 136894
rect 495502 136658 495586 136894
rect 495822 136658 531266 136894
rect 531502 136658 531586 136894
rect 531822 136658 567266 136894
rect 567502 136658 567586 136894
rect 567822 136658 590142 136894
rect 590378 136658 590462 136894
rect 590698 136658 590730 136894
rect -6806 136574 590730 136658
rect -6806 136338 -6774 136574
rect -6538 136338 -6454 136574
rect -6218 136338 27266 136574
rect 27502 136338 27586 136574
rect 27822 136338 63266 136574
rect 63502 136338 63586 136574
rect 63822 136338 99266 136574
rect 99502 136338 99586 136574
rect 99822 136338 135266 136574
rect 135502 136338 135586 136574
rect 135822 136338 171266 136574
rect 171502 136338 171586 136574
rect 171822 136338 207266 136574
rect 207502 136338 207586 136574
rect 207822 136338 243266 136574
rect 243502 136338 243586 136574
rect 243822 136338 279266 136574
rect 279502 136338 279586 136574
rect 279822 136338 315266 136574
rect 315502 136338 315586 136574
rect 315822 136338 351266 136574
rect 351502 136338 351586 136574
rect 351822 136338 387266 136574
rect 387502 136338 387586 136574
rect 387822 136338 423266 136574
rect 423502 136338 423586 136574
rect 423822 136338 459266 136574
rect 459502 136338 459586 136574
rect 459822 136338 495266 136574
rect 495502 136338 495586 136574
rect 495822 136338 531266 136574
rect 531502 136338 531586 136574
rect 531822 136338 567266 136574
rect 567502 136338 567586 136574
rect 567822 136338 590142 136574
rect 590378 136338 590462 136574
rect 590698 136338 590730 136574
rect -6806 136306 590730 136338
rect -4886 133174 588810 133206
rect -4886 132938 -4854 133174
rect -4618 132938 -4534 133174
rect -4298 132938 23546 133174
rect 23782 132938 23866 133174
rect 24102 132938 59546 133174
rect 59782 132938 59866 133174
rect 60102 132938 95546 133174
rect 95782 132938 95866 133174
rect 96102 132938 131546 133174
rect 131782 132938 131866 133174
rect 132102 132938 167546 133174
rect 167782 132938 167866 133174
rect 168102 132938 203546 133174
rect 203782 132938 203866 133174
rect 204102 132938 239546 133174
rect 239782 132938 239866 133174
rect 240102 132938 275546 133174
rect 275782 132938 275866 133174
rect 276102 132938 311546 133174
rect 311782 132938 311866 133174
rect 312102 132938 347546 133174
rect 347782 132938 347866 133174
rect 348102 132938 383546 133174
rect 383782 132938 383866 133174
rect 384102 132938 419546 133174
rect 419782 132938 419866 133174
rect 420102 132938 455546 133174
rect 455782 132938 455866 133174
rect 456102 132938 491546 133174
rect 491782 132938 491866 133174
rect 492102 132938 527546 133174
rect 527782 132938 527866 133174
rect 528102 132938 563546 133174
rect 563782 132938 563866 133174
rect 564102 132938 588222 133174
rect 588458 132938 588542 133174
rect 588778 132938 588810 133174
rect -4886 132854 588810 132938
rect -4886 132618 -4854 132854
rect -4618 132618 -4534 132854
rect -4298 132618 23546 132854
rect 23782 132618 23866 132854
rect 24102 132618 59546 132854
rect 59782 132618 59866 132854
rect 60102 132618 95546 132854
rect 95782 132618 95866 132854
rect 96102 132618 131546 132854
rect 131782 132618 131866 132854
rect 132102 132618 167546 132854
rect 167782 132618 167866 132854
rect 168102 132618 203546 132854
rect 203782 132618 203866 132854
rect 204102 132618 239546 132854
rect 239782 132618 239866 132854
rect 240102 132618 275546 132854
rect 275782 132618 275866 132854
rect 276102 132618 311546 132854
rect 311782 132618 311866 132854
rect 312102 132618 347546 132854
rect 347782 132618 347866 132854
rect 348102 132618 383546 132854
rect 383782 132618 383866 132854
rect 384102 132618 419546 132854
rect 419782 132618 419866 132854
rect 420102 132618 455546 132854
rect 455782 132618 455866 132854
rect 456102 132618 491546 132854
rect 491782 132618 491866 132854
rect 492102 132618 527546 132854
rect 527782 132618 527866 132854
rect 528102 132618 563546 132854
rect 563782 132618 563866 132854
rect 564102 132618 588222 132854
rect 588458 132618 588542 132854
rect 588778 132618 588810 132854
rect -4886 132586 588810 132618
rect -2966 129454 586890 129486
rect -2966 129218 -2934 129454
rect -2698 129218 -2614 129454
rect -2378 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 91826 129454
rect 92062 129218 92146 129454
rect 92382 129218 127826 129454
rect 128062 129218 128146 129454
rect 128382 129218 163826 129454
rect 164062 129218 164146 129454
rect 164382 129218 199826 129454
rect 200062 129218 200146 129454
rect 200382 129218 235826 129454
rect 236062 129218 236146 129454
rect 236382 129218 271826 129454
rect 272062 129218 272146 129454
rect 272382 129218 307826 129454
rect 308062 129218 308146 129454
rect 308382 129218 343826 129454
rect 344062 129218 344146 129454
rect 344382 129218 379826 129454
rect 380062 129218 380146 129454
rect 380382 129218 415826 129454
rect 416062 129218 416146 129454
rect 416382 129218 451826 129454
rect 452062 129218 452146 129454
rect 452382 129218 487826 129454
rect 488062 129218 488146 129454
rect 488382 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 586302 129454
rect 586538 129218 586622 129454
rect 586858 129218 586890 129454
rect -2966 129134 586890 129218
rect -2966 128898 -2934 129134
rect -2698 128898 -2614 129134
rect -2378 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 91826 129134
rect 92062 128898 92146 129134
rect 92382 128898 127826 129134
rect 128062 128898 128146 129134
rect 128382 128898 163826 129134
rect 164062 128898 164146 129134
rect 164382 128898 199826 129134
rect 200062 128898 200146 129134
rect 200382 128898 235826 129134
rect 236062 128898 236146 129134
rect 236382 128898 271826 129134
rect 272062 128898 272146 129134
rect 272382 128898 307826 129134
rect 308062 128898 308146 129134
rect 308382 128898 343826 129134
rect 344062 128898 344146 129134
rect 344382 128898 379826 129134
rect 380062 128898 380146 129134
rect 380382 128898 415826 129134
rect 416062 128898 416146 129134
rect 416382 128898 451826 129134
rect 452062 128898 452146 129134
rect 452382 128898 487826 129134
rect 488062 128898 488146 129134
rect 488382 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 586302 129134
rect 586538 128898 586622 129134
rect 586858 128898 586890 129134
rect -2966 128866 586890 128898
rect -8726 122614 592650 122646
rect -8726 122378 -7734 122614
rect -7498 122378 -7414 122614
rect -7178 122378 12986 122614
rect 13222 122378 13306 122614
rect 13542 122378 48986 122614
rect 49222 122378 49306 122614
rect 49542 122378 84986 122614
rect 85222 122378 85306 122614
rect 85542 122378 120986 122614
rect 121222 122378 121306 122614
rect 121542 122378 156986 122614
rect 157222 122378 157306 122614
rect 157542 122378 192986 122614
rect 193222 122378 193306 122614
rect 193542 122378 228986 122614
rect 229222 122378 229306 122614
rect 229542 122378 264986 122614
rect 265222 122378 265306 122614
rect 265542 122378 300986 122614
rect 301222 122378 301306 122614
rect 301542 122378 336986 122614
rect 337222 122378 337306 122614
rect 337542 122378 372986 122614
rect 373222 122378 373306 122614
rect 373542 122378 408986 122614
rect 409222 122378 409306 122614
rect 409542 122378 444986 122614
rect 445222 122378 445306 122614
rect 445542 122378 480986 122614
rect 481222 122378 481306 122614
rect 481542 122378 516986 122614
rect 517222 122378 517306 122614
rect 517542 122378 552986 122614
rect 553222 122378 553306 122614
rect 553542 122378 591102 122614
rect 591338 122378 591422 122614
rect 591658 122378 592650 122614
rect -8726 122294 592650 122378
rect -8726 122058 -7734 122294
rect -7498 122058 -7414 122294
rect -7178 122058 12986 122294
rect 13222 122058 13306 122294
rect 13542 122058 48986 122294
rect 49222 122058 49306 122294
rect 49542 122058 84986 122294
rect 85222 122058 85306 122294
rect 85542 122058 120986 122294
rect 121222 122058 121306 122294
rect 121542 122058 156986 122294
rect 157222 122058 157306 122294
rect 157542 122058 192986 122294
rect 193222 122058 193306 122294
rect 193542 122058 228986 122294
rect 229222 122058 229306 122294
rect 229542 122058 264986 122294
rect 265222 122058 265306 122294
rect 265542 122058 300986 122294
rect 301222 122058 301306 122294
rect 301542 122058 336986 122294
rect 337222 122058 337306 122294
rect 337542 122058 372986 122294
rect 373222 122058 373306 122294
rect 373542 122058 408986 122294
rect 409222 122058 409306 122294
rect 409542 122058 444986 122294
rect 445222 122058 445306 122294
rect 445542 122058 480986 122294
rect 481222 122058 481306 122294
rect 481542 122058 516986 122294
rect 517222 122058 517306 122294
rect 517542 122058 552986 122294
rect 553222 122058 553306 122294
rect 553542 122058 591102 122294
rect 591338 122058 591422 122294
rect 591658 122058 592650 122294
rect -8726 122026 592650 122058
rect -6806 118894 590730 118926
rect -6806 118658 -5814 118894
rect -5578 118658 -5494 118894
rect -5258 118658 9266 118894
rect 9502 118658 9586 118894
rect 9822 118658 45266 118894
rect 45502 118658 45586 118894
rect 45822 118658 81266 118894
rect 81502 118658 81586 118894
rect 81822 118658 117266 118894
rect 117502 118658 117586 118894
rect 117822 118658 153266 118894
rect 153502 118658 153586 118894
rect 153822 118658 189266 118894
rect 189502 118658 189586 118894
rect 189822 118658 225266 118894
rect 225502 118658 225586 118894
rect 225822 118658 261266 118894
rect 261502 118658 261586 118894
rect 261822 118658 297266 118894
rect 297502 118658 297586 118894
rect 297822 118658 333266 118894
rect 333502 118658 333586 118894
rect 333822 118658 369266 118894
rect 369502 118658 369586 118894
rect 369822 118658 405266 118894
rect 405502 118658 405586 118894
rect 405822 118658 441266 118894
rect 441502 118658 441586 118894
rect 441822 118658 477266 118894
rect 477502 118658 477586 118894
rect 477822 118658 513266 118894
rect 513502 118658 513586 118894
rect 513822 118658 549266 118894
rect 549502 118658 549586 118894
rect 549822 118658 589182 118894
rect 589418 118658 589502 118894
rect 589738 118658 590730 118894
rect -6806 118574 590730 118658
rect -6806 118338 -5814 118574
rect -5578 118338 -5494 118574
rect -5258 118338 9266 118574
rect 9502 118338 9586 118574
rect 9822 118338 45266 118574
rect 45502 118338 45586 118574
rect 45822 118338 81266 118574
rect 81502 118338 81586 118574
rect 81822 118338 117266 118574
rect 117502 118338 117586 118574
rect 117822 118338 153266 118574
rect 153502 118338 153586 118574
rect 153822 118338 189266 118574
rect 189502 118338 189586 118574
rect 189822 118338 225266 118574
rect 225502 118338 225586 118574
rect 225822 118338 261266 118574
rect 261502 118338 261586 118574
rect 261822 118338 297266 118574
rect 297502 118338 297586 118574
rect 297822 118338 333266 118574
rect 333502 118338 333586 118574
rect 333822 118338 369266 118574
rect 369502 118338 369586 118574
rect 369822 118338 405266 118574
rect 405502 118338 405586 118574
rect 405822 118338 441266 118574
rect 441502 118338 441586 118574
rect 441822 118338 477266 118574
rect 477502 118338 477586 118574
rect 477822 118338 513266 118574
rect 513502 118338 513586 118574
rect 513822 118338 549266 118574
rect 549502 118338 549586 118574
rect 549822 118338 589182 118574
rect 589418 118338 589502 118574
rect 589738 118338 590730 118574
rect -6806 118306 590730 118338
rect -4886 115174 588810 115206
rect -4886 114938 -3894 115174
rect -3658 114938 -3574 115174
rect -3338 114938 5546 115174
rect 5782 114938 5866 115174
rect 6102 114938 41546 115174
rect 41782 114938 41866 115174
rect 42102 114938 77546 115174
rect 77782 114938 77866 115174
rect 78102 114938 113546 115174
rect 113782 114938 113866 115174
rect 114102 114938 149546 115174
rect 149782 114938 149866 115174
rect 150102 114938 185546 115174
rect 185782 114938 185866 115174
rect 186102 114938 221546 115174
rect 221782 114938 221866 115174
rect 222102 114938 257546 115174
rect 257782 114938 257866 115174
rect 258102 114938 293546 115174
rect 293782 114938 293866 115174
rect 294102 114938 329546 115174
rect 329782 114938 329866 115174
rect 330102 114938 365546 115174
rect 365782 114938 365866 115174
rect 366102 114938 401546 115174
rect 401782 114938 401866 115174
rect 402102 114938 437546 115174
rect 437782 114938 437866 115174
rect 438102 114938 473546 115174
rect 473782 114938 473866 115174
rect 474102 114938 509546 115174
rect 509782 114938 509866 115174
rect 510102 114938 545546 115174
rect 545782 114938 545866 115174
rect 546102 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 587262 115174
rect 587498 114938 587582 115174
rect 587818 114938 588810 115174
rect -4886 114854 588810 114938
rect -4886 114618 -3894 114854
rect -3658 114618 -3574 114854
rect -3338 114618 5546 114854
rect 5782 114618 5866 114854
rect 6102 114618 41546 114854
rect 41782 114618 41866 114854
rect 42102 114618 77546 114854
rect 77782 114618 77866 114854
rect 78102 114618 113546 114854
rect 113782 114618 113866 114854
rect 114102 114618 149546 114854
rect 149782 114618 149866 114854
rect 150102 114618 185546 114854
rect 185782 114618 185866 114854
rect 186102 114618 221546 114854
rect 221782 114618 221866 114854
rect 222102 114618 257546 114854
rect 257782 114618 257866 114854
rect 258102 114618 293546 114854
rect 293782 114618 293866 114854
rect 294102 114618 329546 114854
rect 329782 114618 329866 114854
rect 330102 114618 365546 114854
rect 365782 114618 365866 114854
rect 366102 114618 401546 114854
rect 401782 114618 401866 114854
rect 402102 114618 437546 114854
rect 437782 114618 437866 114854
rect 438102 114618 473546 114854
rect 473782 114618 473866 114854
rect 474102 114618 509546 114854
rect 509782 114618 509866 114854
rect 510102 114618 545546 114854
rect 545782 114618 545866 114854
rect 546102 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 587262 114854
rect 587498 114618 587582 114854
rect 587818 114618 588810 114854
rect -4886 114586 588810 114618
rect -2966 111454 586890 111486
rect -2966 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 73826 111454
rect 74062 111218 74146 111454
rect 74382 111218 109826 111454
rect 110062 111218 110146 111454
rect 110382 111218 145826 111454
rect 146062 111218 146146 111454
rect 146382 111218 181826 111454
rect 182062 111218 182146 111454
rect 182382 111218 217826 111454
rect 218062 111218 218146 111454
rect 218382 111218 253826 111454
rect 254062 111218 254146 111454
rect 254382 111218 289826 111454
rect 290062 111218 290146 111454
rect 290382 111218 325826 111454
rect 326062 111218 326146 111454
rect 326382 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 586890 111454
rect -2966 111134 586890 111218
rect -2966 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 73826 111134
rect 74062 110898 74146 111134
rect 74382 110898 109826 111134
rect 110062 110898 110146 111134
rect 110382 110898 145826 111134
rect 146062 110898 146146 111134
rect 146382 110898 181826 111134
rect 182062 110898 182146 111134
rect 182382 110898 217826 111134
rect 218062 110898 218146 111134
rect 218382 110898 253826 111134
rect 254062 110898 254146 111134
rect 254382 110898 289826 111134
rect 290062 110898 290146 111134
rect 290382 110898 325826 111134
rect 326062 110898 326146 111134
rect 326382 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 586890 111134
rect -2966 110866 586890 110898
rect -8726 104614 592650 104646
rect -8726 104378 -8694 104614
rect -8458 104378 -8374 104614
rect -8138 104378 30986 104614
rect 31222 104378 31306 104614
rect 31542 104378 66986 104614
rect 67222 104378 67306 104614
rect 67542 104378 102986 104614
rect 103222 104378 103306 104614
rect 103542 104378 138986 104614
rect 139222 104378 139306 104614
rect 139542 104378 174986 104614
rect 175222 104378 175306 104614
rect 175542 104378 210986 104614
rect 211222 104378 211306 104614
rect 211542 104378 246986 104614
rect 247222 104378 247306 104614
rect 247542 104378 282986 104614
rect 283222 104378 283306 104614
rect 283542 104378 318986 104614
rect 319222 104378 319306 104614
rect 319542 104378 354986 104614
rect 355222 104378 355306 104614
rect 355542 104378 390986 104614
rect 391222 104378 391306 104614
rect 391542 104378 426986 104614
rect 427222 104378 427306 104614
rect 427542 104378 462986 104614
rect 463222 104378 463306 104614
rect 463542 104378 498986 104614
rect 499222 104378 499306 104614
rect 499542 104378 534986 104614
rect 535222 104378 535306 104614
rect 535542 104378 570986 104614
rect 571222 104378 571306 104614
rect 571542 104378 592062 104614
rect 592298 104378 592382 104614
rect 592618 104378 592650 104614
rect -8726 104294 592650 104378
rect -8726 104058 -8694 104294
rect -8458 104058 -8374 104294
rect -8138 104058 30986 104294
rect 31222 104058 31306 104294
rect 31542 104058 66986 104294
rect 67222 104058 67306 104294
rect 67542 104058 102986 104294
rect 103222 104058 103306 104294
rect 103542 104058 138986 104294
rect 139222 104058 139306 104294
rect 139542 104058 174986 104294
rect 175222 104058 175306 104294
rect 175542 104058 210986 104294
rect 211222 104058 211306 104294
rect 211542 104058 246986 104294
rect 247222 104058 247306 104294
rect 247542 104058 282986 104294
rect 283222 104058 283306 104294
rect 283542 104058 318986 104294
rect 319222 104058 319306 104294
rect 319542 104058 354986 104294
rect 355222 104058 355306 104294
rect 355542 104058 390986 104294
rect 391222 104058 391306 104294
rect 391542 104058 426986 104294
rect 427222 104058 427306 104294
rect 427542 104058 462986 104294
rect 463222 104058 463306 104294
rect 463542 104058 498986 104294
rect 499222 104058 499306 104294
rect 499542 104058 534986 104294
rect 535222 104058 535306 104294
rect 535542 104058 570986 104294
rect 571222 104058 571306 104294
rect 571542 104058 592062 104294
rect 592298 104058 592382 104294
rect 592618 104058 592650 104294
rect -8726 104026 592650 104058
rect -6806 100894 590730 100926
rect -6806 100658 -6774 100894
rect -6538 100658 -6454 100894
rect -6218 100658 27266 100894
rect 27502 100658 27586 100894
rect 27822 100658 63266 100894
rect 63502 100658 63586 100894
rect 63822 100658 99266 100894
rect 99502 100658 99586 100894
rect 99822 100658 135266 100894
rect 135502 100658 135586 100894
rect 135822 100658 171266 100894
rect 171502 100658 171586 100894
rect 171822 100658 207266 100894
rect 207502 100658 207586 100894
rect 207822 100658 243266 100894
rect 243502 100658 243586 100894
rect 243822 100658 279266 100894
rect 279502 100658 279586 100894
rect 279822 100658 315266 100894
rect 315502 100658 315586 100894
rect 315822 100658 351266 100894
rect 351502 100658 351586 100894
rect 351822 100658 387266 100894
rect 387502 100658 387586 100894
rect 387822 100658 423266 100894
rect 423502 100658 423586 100894
rect 423822 100658 459266 100894
rect 459502 100658 459586 100894
rect 459822 100658 495266 100894
rect 495502 100658 495586 100894
rect 495822 100658 531266 100894
rect 531502 100658 531586 100894
rect 531822 100658 567266 100894
rect 567502 100658 567586 100894
rect 567822 100658 590142 100894
rect 590378 100658 590462 100894
rect 590698 100658 590730 100894
rect -6806 100574 590730 100658
rect -6806 100338 -6774 100574
rect -6538 100338 -6454 100574
rect -6218 100338 27266 100574
rect 27502 100338 27586 100574
rect 27822 100338 63266 100574
rect 63502 100338 63586 100574
rect 63822 100338 99266 100574
rect 99502 100338 99586 100574
rect 99822 100338 135266 100574
rect 135502 100338 135586 100574
rect 135822 100338 171266 100574
rect 171502 100338 171586 100574
rect 171822 100338 207266 100574
rect 207502 100338 207586 100574
rect 207822 100338 243266 100574
rect 243502 100338 243586 100574
rect 243822 100338 279266 100574
rect 279502 100338 279586 100574
rect 279822 100338 315266 100574
rect 315502 100338 315586 100574
rect 315822 100338 351266 100574
rect 351502 100338 351586 100574
rect 351822 100338 387266 100574
rect 387502 100338 387586 100574
rect 387822 100338 423266 100574
rect 423502 100338 423586 100574
rect 423822 100338 459266 100574
rect 459502 100338 459586 100574
rect 459822 100338 495266 100574
rect 495502 100338 495586 100574
rect 495822 100338 531266 100574
rect 531502 100338 531586 100574
rect 531822 100338 567266 100574
rect 567502 100338 567586 100574
rect 567822 100338 590142 100574
rect 590378 100338 590462 100574
rect 590698 100338 590730 100574
rect -6806 100306 590730 100338
rect -4886 97174 588810 97206
rect -4886 96938 -4854 97174
rect -4618 96938 -4534 97174
rect -4298 96938 23546 97174
rect 23782 96938 23866 97174
rect 24102 96938 59546 97174
rect 59782 96938 59866 97174
rect 60102 96938 95546 97174
rect 95782 96938 95866 97174
rect 96102 96938 131546 97174
rect 131782 96938 131866 97174
rect 132102 96938 167546 97174
rect 167782 96938 167866 97174
rect 168102 96938 203546 97174
rect 203782 96938 203866 97174
rect 204102 96938 239546 97174
rect 239782 96938 239866 97174
rect 240102 96938 275546 97174
rect 275782 96938 275866 97174
rect 276102 96938 311546 97174
rect 311782 96938 311866 97174
rect 312102 96938 347546 97174
rect 347782 96938 347866 97174
rect 348102 96938 383546 97174
rect 383782 96938 383866 97174
rect 384102 96938 419546 97174
rect 419782 96938 419866 97174
rect 420102 96938 455546 97174
rect 455782 96938 455866 97174
rect 456102 96938 491546 97174
rect 491782 96938 491866 97174
rect 492102 96938 527546 97174
rect 527782 96938 527866 97174
rect 528102 96938 563546 97174
rect 563782 96938 563866 97174
rect 564102 96938 588222 97174
rect 588458 96938 588542 97174
rect 588778 96938 588810 97174
rect -4886 96854 588810 96938
rect -4886 96618 -4854 96854
rect -4618 96618 -4534 96854
rect -4298 96618 23546 96854
rect 23782 96618 23866 96854
rect 24102 96618 59546 96854
rect 59782 96618 59866 96854
rect 60102 96618 95546 96854
rect 95782 96618 95866 96854
rect 96102 96618 131546 96854
rect 131782 96618 131866 96854
rect 132102 96618 167546 96854
rect 167782 96618 167866 96854
rect 168102 96618 203546 96854
rect 203782 96618 203866 96854
rect 204102 96618 239546 96854
rect 239782 96618 239866 96854
rect 240102 96618 275546 96854
rect 275782 96618 275866 96854
rect 276102 96618 311546 96854
rect 311782 96618 311866 96854
rect 312102 96618 347546 96854
rect 347782 96618 347866 96854
rect 348102 96618 383546 96854
rect 383782 96618 383866 96854
rect 384102 96618 419546 96854
rect 419782 96618 419866 96854
rect 420102 96618 455546 96854
rect 455782 96618 455866 96854
rect 456102 96618 491546 96854
rect 491782 96618 491866 96854
rect 492102 96618 527546 96854
rect 527782 96618 527866 96854
rect 528102 96618 563546 96854
rect 563782 96618 563866 96854
rect 564102 96618 588222 96854
rect 588458 96618 588542 96854
rect 588778 96618 588810 96854
rect -4886 96586 588810 96618
rect -2966 93454 586890 93486
rect -2966 93218 -2934 93454
rect -2698 93218 -2614 93454
rect -2378 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 91826 93454
rect 92062 93218 92146 93454
rect 92382 93218 127826 93454
rect 128062 93218 128146 93454
rect 128382 93218 163826 93454
rect 164062 93218 164146 93454
rect 164382 93218 199826 93454
rect 200062 93218 200146 93454
rect 200382 93218 235826 93454
rect 236062 93218 236146 93454
rect 236382 93218 271826 93454
rect 272062 93218 272146 93454
rect 272382 93218 307826 93454
rect 308062 93218 308146 93454
rect 308382 93218 343826 93454
rect 344062 93218 344146 93454
rect 344382 93218 379826 93454
rect 380062 93218 380146 93454
rect 380382 93218 415826 93454
rect 416062 93218 416146 93454
rect 416382 93218 451826 93454
rect 452062 93218 452146 93454
rect 452382 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 586302 93454
rect 586538 93218 586622 93454
rect 586858 93218 586890 93454
rect -2966 93134 586890 93218
rect -2966 92898 -2934 93134
rect -2698 92898 -2614 93134
rect -2378 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 91826 93134
rect 92062 92898 92146 93134
rect 92382 92898 127826 93134
rect 128062 92898 128146 93134
rect 128382 92898 163826 93134
rect 164062 92898 164146 93134
rect 164382 92898 199826 93134
rect 200062 92898 200146 93134
rect 200382 92898 235826 93134
rect 236062 92898 236146 93134
rect 236382 92898 271826 93134
rect 272062 92898 272146 93134
rect 272382 92898 307826 93134
rect 308062 92898 308146 93134
rect 308382 92898 343826 93134
rect 344062 92898 344146 93134
rect 344382 92898 379826 93134
rect 380062 92898 380146 93134
rect 380382 92898 415826 93134
rect 416062 92898 416146 93134
rect 416382 92898 451826 93134
rect 452062 92898 452146 93134
rect 452382 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 586302 93134
rect 586538 92898 586622 93134
rect 586858 92898 586890 93134
rect -2966 92866 586890 92898
rect -8726 86614 592650 86646
rect -8726 86378 -7734 86614
rect -7498 86378 -7414 86614
rect -7178 86378 12986 86614
rect 13222 86378 13306 86614
rect 13542 86378 48986 86614
rect 49222 86378 49306 86614
rect 49542 86378 84986 86614
rect 85222 86378 85306 86614
rect 85542 86378 120986 86614
rect 121222 86378 121306 86614
rect 121542 86378 156986 86614
rect 157222 86378 157306 86614
rect 157542 86378 192986 86614
rect 193222 86378 193306 86614
rect 193542 86378 228986 86614
rect 229222 86378 229306 86614
rect 229542 86378 264986 86614
rect 265222 86378 265306 86614
rect 265542 86378 300986 86614
rect 301222 86378 301306 86614
rect 301542 86378 336986 86614
rect 337222 86378 337306 86614
rect 337542 86378 372986 86614
rect 373222 86378 373306 86614
rect 373542 86378 408986 86614
rect 409222 86378 409306 86614
rect 409542 86378 444986 86614
rect 445222 86378 445306 86614
rect 445542 86378 480986 86614
rect 481222 86378 481306 86614
rect 481542 86378 516986 86614
rect 517222 86378 517306 86614
rect 517542 86378 552986 86614
rect 553222 86378 553306 86614
rect 553542 86378 591102 86614
rect 591338 86378 591422 86614
rect 591658 86378 592650 86614
rect -8726 86294 592650 86378
rect -8726 86058 -7734 86294
rect -7498 86058 -7414 86294
rect -7178 86058 12986 86294
rect 13222 86058 13306 86294
rect 13542 86058 48986 86294
rect 49222 86058 49306 86294
rect 49542 86058 84986 86294
rect 85222 86058 85306 86294
rect 85542 86058 120986 86294
rect 121222 86058 121306 86294
rect 121542 86058 156986 86294
rect 157222 86058 157306 86294
rect 157542 86058 192986 86294
rect 193222 86058 193306 86294
rect 193542 86058 228986 86294
rect 229222 86058 229306 86294
rect 229542 86058 264986 86294
rect 265222 86058 265306 86294
rect 265542 86058 300986 86294
rect 301222 86058 301306 86294
rect 301542 86058 336986 86294
rect 337222 86058 337306 86294
rect 337542 86058 372986 86294
rect 373222 86058 373306 86294
rect 373542 86058 408986 86294
rect 409222 86058 409306 86294
rect 409542 86058 444986 86294
rect 445222 86058 445306 86294
rect 445542 86058 480986 86294
rect 481222 86058 481306 86294
rect 481542 86058 516986 86294
rect 517222 86058 517306 86294
rect 517542 86058 552986 86294
rect 553222 86058 553306 86294
rect 553542 86058 591102 86294
rect 591338 86058 591422 86294
rect 591658 86058 592650 86294
rect -8726 86026 592650 86058
rect -6806 82894 590730 82926
rect -6806 82658 -5814 82894
rect -5578 82658 -5494 82894
rect -5258 82658 9266 82894
rect 9502 82658 9586 82894
rect 9822 82658 45266 82894
rect 45502 82658 45586 82894
rect 45822 82658 81266 82894
rect 81502 82658 81586 82894
rect 81822 82658 117266 82894
rect 117502 82658 117586 82894
rect 117822 82658 153266 82894
rect 153502 82658 153586 82894
rect 153822 82658 189266 82894
rect 189502 82658 189586 82894
rect 189822 82658 225266 82894
rect 225502 82658 225586 82894
rect 225822 82658 261266 82894
rect 261502 82658 261586 82894
rect 261822 82658 297266 82894
rect 297502 82658 297586 82894
rect 297822 82658 333266 82894
rect 333502 82658 333586 82894
rect 333822 82658 369266 82894
rect 369502 82658 369586 82894
rect 369822 82658 405266 82894
rect 405502 82658 405586 82894
rect 405822 82658 441266 82894
rect 441502 82658 441586 82894
rect 441822 82658 477266 82894
rect 477502 82658 477586 82894
rect 477822 82658 513266 82894
rect 513502 82658 513586 82894
rect 513822 82658 549266 82894
rect 549502 82658 549586 82894
rect 549822 82658 589182 82894
rect 589418 82658 589502 82894
rect 589738 82658 590730 82894
rect -6806 82574 590730 82658
rect -6806 82338 -5814 82574
rect -5578 82338 -5494 82574
rect -5258 82338 9266 82574
rect 9502 82338 9586 82574
rect 9822 82338 45266 82574
rect 45502 82338 45586 82574
rect 45822 82338 81266 82574
rect 81502 82338 81586 82574
rect 81822 82338 117266 82574
rect 117502 82338 117586 82574
rect 117822 82338 153266 82574
rect 153502 82338 153586 82574
rect 153822 82338 189266 82574
rect 189502 82338 189586 82574
rect 189822 82338 225266 82574
rect 225502 82338 225586 82574
rect 225822 82338 261266 82574
rect 261502 82338 261586 82574
rect 261822 82338 297266 82574
rect 297502 82338 297586 82574
rect 297822 82338 333266 82574
rect 333502 82338 333586 82574
rect 333822 82338 369266 82574
rect 369502 82338 369586 82574
rect 369822 82338 405266 82574
rect 405502 82338 405586 82574
rect 405822 82338 441266 82574
rect 441502 82338 441586 82574
rect 441822 82338 477266 82574
rect 477502 82338 477586 82574
rect 477822 82338 513266 82574
rect 513502 82338 513586 82574
rect 513822 82338 549266 82574
rect 549502 82338 549586 82574
rect 549822 82338 589182 82574
rect 589418 82338 589502 82574
rect 589738 82338 590730 82574
rect -6806 82306 590730 82338
rect -4886 79174 588810 79206
rect -4886 78938 -3894 79174
rect -3658 78938 -3574 79174
rect -3338 78938 5546 79174
rect 5782 78938 5866 79174
rect 6102 78938 41546 79174
rect 41782 78938 41866 79174
rect 42102 78938 77546 79174
rect 77782 78938 77866 79174
rect 78102 78938 113546 79174
rect 113782 78938 113866 79174
rect 114102 78938 149546 79174
rect 149782 78938 149866 79174
rect 150102 78938 185546 79174
rect 185782 78938 185866 79174
rect 186102 78938 221546 79174
rect 221782 78938 221866 79174
rect 222102 78938 257546 79174
rect 257782 78938 257866 79174
rect 258102 78938 293546 79174
rect 293782 78938 293866 79174
rect 294102 78938 329546 79174
rect 329782 78938 329866 79174
rect 330102 78938 365546 79174
rect 365782 78938 365866 79174
rect 366102 78938 401546 79174
rect 401782 78938 401866 79174
rect 402102 78938 437546 79174
rect 437782 78938 437866 79174
rect 438102 78938 473546 79174
rect 473782 78938 473866 79174
rect 474102 78938 509546 79174
rect 509782 78938 509866 79174
rect 510102 78938 545546 79174
rect 545782 78938 545866 79174
rect 546102 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 587262 79174
rect 587498 78938 587582 79174
rect 587818 78938 588810 79174
rect -4886 78854 588810 78938
rect -4886 78618 -3894 78854
rect -3658 78618 -3574 78854
rect -3338 78618 5546 78854
rect 5782 78618 5866 78854
rect 6102 78618 41546 78854
rect 41782 78618 41866 78854
rect 42102 78618 77546 78854
rect 77782 78618 77866 78854
rect 78102 78618 113546 78854
rect 113782 78618 113866 78854
rect 114102 78618 149546 78854
rect 149782 78618 149866 78854
rect 150102 78618 185546 78854
rect 185782 78618 185866 78854
rect 186102 78618 221546 78854
rect 221782 78618 221866 78854
rect 222102 78618 257546 78854
rect 257782 78618 257866 78854
rect 258102 78618 293546 78854
rect 293782 78618 293866 78854
rect 294102 78618 329546 78854
rect 329782 78618 329866 78854
rect 330102 78618 365546 78854
rect 365782 78618 365866 78854
rect 366102 78618 401546 78854
rect 401782 78618 401866 78854
rect 402102 78618 437546 78854
rect 437782 78618 437866 78854
rect 438102 78618 473546 78854
rect 473782 78618 473866 78854
rect 474102 78618 509546 78854
rect 509782 78618 509866 78854
rect 510102 78618 545546 78854
rect 545782 78618 545866 78854
rect 546102 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 587262 78854
rect 587498 78618 587582 78854
rect 587818 78618 588810 78854
rect -4886 78586 588810 78618
rect -2966 75454 586890 75486
rect -2966 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 73826 75454
rect 74062 75218 74146 75454
rect 74382 75218 109826 75454
rect 110062 75218 110146 75454
rect 110382 75218 145826 75454
rect 146062 75218 146146 75454
rect 146382 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 217826 75454
rect 218062 75218 218146 75454
rect 218382 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 586890 75454
rect -2966 75134 586890 75218
rect -2966 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 73826 75134
rect 74062 74898 74146 75134
rect 74382 74898 109826 75134
rect 110062 74898 110146 75134
rect 110382 74898 145826 75134
rect 146062 74898 146146 75134
rect 146382 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 217826 75134
rect 218062 74898 218146 75134
rect 218382 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 586890 75134
rect -2966 74866 586890 74898
rect -8726 68614 592650 68646
rect -8726 68378 -8694 68614
rect -8458 68378 -8374 68614
rect -8138 68378 30986 68614
rect 31222 68378 31306 68614
rect 31542 68378 66986 68614
rect 67222 68378 67306 68614
rect 67542 68378 102986 68614
rect 103222 68378 103306 68614
rect 103542 68378 138986 68614
rect 139222 68378 139306 68614
rect 139542 68378 174986 68614
rect 175222 68378 175306 68614
rect 175542 68378 210986 68614
rect 211222 68378 211306 68614
rect 211542 68378 246986 68614
rect 247222 68378 247306 68614
rect 247542 68378 282986 68614
rect 283222 68378 283306 68614
rect 283542 68378 318986 68614
rect 319222 68378 319306 68614
rect 319542 68378 354986 68614
rect 355222 68378 355306 68614
rect 355542 68378 390986 68614
rect 391222 68378 391306 68614
rect 391542 68378 426986 68614
rect 427222 68378 427306 68614
rect 427542 68378 462986 68614
rect 463222 68378 463306 68614
rect 463542 68378 498986 68614
rect 499222 68378 499306 68614
rect 499542 68378 534986 68614
rect 535222 68378 535306 68614
rect 535542 68378 570986 68614
rect 571222 68378 571306 68614
rect 571542 68378 592062 68614
rect 592298 68378 592382 68614
rect 592618 68378 592650 68614
rect -8726 68294 592650 68378
rect -8726 68058 -8694 68294
rect -8458 68058 -8374 68294
rect -8138 68058 30986 68294
rect 31222 68058 31306 68294
rect 31542 68058 66986 68294
rect 67222 68058 67306 68294
rect 67542 68058 102986 68294
rect 103222 68058 103306 68294
rect 103542 68058 138986 68294
rect 139222 68058 139306 68294
rect 139542 68058 174986 68294
rect 175222 68058 175306 68294
rect 175542 68058 210986 68294
rect 211222 68058 211306 68294
rect 211542 68058 246986 68294
rect 247222 68058 247306 68294
rect 247542 68058 282986 68294
rect 283222 68058 283306 68294
rect 283542 68058 318986 68294
rect 319222 68058 319306 68294
rect 319542 68058 354986 68294
rect 355222 68058 355306 68294
rect 355542 68058 390986 68294
rect 391222 68058 391306 68294
rect 391542 68058 426986 68294
rect 427222 68058 427306 68294
rect 427542 68058 462986 68294
rect 463222 68058 463306 68294
rect 463542 68058 498986 68294
rect 499222 68058 499306 68294
rect 499542 68058 534986 68294
rect 535222 68058 535306 68294
rect 535542 68058 570986 68294
rect 571222 68058 571306 68294
rect 571542 68058 592062 68294
rect 592298 68058 592382 68294
rect 592618 68058 592650 68294
rect -8726 68026 592650 68058
rect -6806 64894 590730 64926
rect -6806 64658 -6774 64894
rect -6538 64658 -6454 64894
rect -6218 64658 27266 64894
rect 27502 64658 27586 64894
rect 27822 64658 63266 64894
rect 63502 64658 63586 64894
rect 63822 64658 99266 64894
rect 99502 64658 99586 64894
rect 99822 64658 135266 64894
rect 135502 64658 135586 64894
rect 135822 64658 171266 64894
rect 171502 64658 171586 64894
rect 171822 64658 207266 64894
rect 207502 64658 207586 64894
rect 207822 64658 243266 64894
rect 243502 64658 243586 64894
rect 243822 64658 279266 64894
rect 279502 64658 279586 64894
rect 279822 64658 315266 64894
rect 315502 64658 315586 64894
rect 315822 64658 351266 64894
rect 351502 64658 351586 64894
rect 351822 64658 387266 64894
rect 387502 64658 387586 64894
rect 387822 64658 423266 64894
rect 423502 64658 423586 64894
rect 423822 64658 459266 64894
rect 459502 64658 459586 64894
rect 459822 64658 495266 64894
rect 495502 64658 495586 64894
rect 495822 64658 531266 64894
rect 531502 64658 531586 64894
rect 531822 64658 567266 64894
rect 567502 64658 567586 64894
rect 567822 64658 590142 64894
rect 590378 64658 590462 64894
rect 590698 64658 590730 64894
rect -6806 64574 590730 64658
rect -6806 64338 -6774 64574
rect -6538 64338 -6454 64574
rect -6218 64338 27266 64574
rect 27502 64338 27586 64574
rect 27822 64338 63266 64574
rect 63502 64338 63586 64574
rect 63822 64338 99266 64574
rect 99502 64338 99586 64574
rect 99822 64338 135266 64574
rect 135502 64338 135586 64574
rect 135822 64338 171266 64574
rect 171502 64338 171586 64574
rect 171822 64338 207266 64574
rect 207502 64338 207586 64574
rect 207822 64338 243266 64574
rect 243502 64338 243586 64574
rect 243822 64338 279266 64574
rect 279502 64338 279586 64574
rect 279822 64338 315266 64574
rect 315502 64338 315586 64574
rect 315822 64338 351266 64574
rect 351502 64338 351586 64574
rect 351822 64338 387266 64574
rect 387502 64338 387586 64574
rect 387822 64338 423266 64574
rect 423502 64338 423586 64574
rect 423822 64338 459266 64574
rect 459502 64338 459586 64574
rect 459822 64338 495266 64574
rect 495502 64338 495586 64574
rect 495822 64338 531266 64574
rect 531502 64338 531586 64574
rect 531822 64338 567266 64574
rect 567502 64338 567586 64574
rect 567822 64338 590142 64574
rect 590378 64338 590462 64574
rect 590698 64338 590730 64574
rect -6806 64306 590730 64338
rect -4886 61174 588810 61206
rect -4886 60938 -4854 61174
rect -4618 60938 -4534 61174
rect -4298 60938 23546 61174
rect 23782 60938 23866 61174
rect 24102 60938 59546 61174
rect 59782 60938 59866 61174
rect 60102 60938 95546 61174
rect 95782 60938 95866 61174
rect 96102 60938 131546 61174
rect 131782 60938 131866 61174
rect 132102 60938 167546 61174
rect 167782 60938 167866 61174
rect 168102 60938 203546 61174
rect 203782 60938 203866 61174
rect 204102 60938 239546 61174
rect 239782 60938 239866 61174
rect 240102 60938 275546 61174
rect 275782 60938 275866 61174
rect 276102 60938 311546 61174
rect 311782 60938 311866 61174
rect 312102 60938 347546 61174
rect 347782 60938 347866 61174
rect 348102 60938 383546 61174
rect 383782 60938 383866 61174
rect 384102 60938 419546 61174
rect 419782 60938 419866 61174
rect 420102 60938 455546 61174
rect 455782 60938 455866 61174
rect 456102 60938 491546 61174
rect 491782 60938 491866 61174
rect 492102 60938 527546 61174
rect 527782 60938 527866 61174
rect 528102 60938 563546 61174
rect 563782 60938 563866 61174
rect 564102 60938 588222 61174
rect 588458 60938 588542 61174
rect 588778 60938 588810 61174
rect -4886 60854 588810 60938
rect -4886 60618 -4854 60854
rect -4618 60618 -4534 60854
rect -4298 60618 23546 60854
rect 23782 60618 23866 60854
rect 24102 60618 59546 60854
rect 59782 60618 59866 60854
rect 60102 60618 95546 60854
rect 95782 60618 95866 60854
rect 96102 60618 131546 60854
rect 131782 60618 131866 60854
rect 132102 60618 167546 60854
rect 167782 60618 167866 60854
rect 168102 60618 203546 60854
rect 203782 60618 203866 60854
rect 204102 60618 239546 60854
rect 239782 60618 239866 60854
rect 240102 60618 275546 60854
rect 275782 60618 275866 60854
rect 276102 60618 311546 60854
rect 311782 60618 311866 60854
rect 312102 60618 347546 60854
rect 347782 60618 347866 60854
rect 348102 60618 383546 60854
rect 383782 60618 383866 60854
rect 384102 60618 419546 60854
rect 419782 60618 419866 60854
rect 420102 60618 455546 60854
rect 455782 60618 455866 60854
rect 456102 60618 491546 60854
rect 491782 60618 491866 60854
rect 492102 60618 527546 60854
rect 527782 60618 527866 60854
rect 528102 60618 563546 60854
rect 563782 60618 563866 60854
rect 564102 60618 588222 60854
rect 588458 60618 588542 60854
rect 588778 60618 588810 60854
rect -4886 60586 588810 60618
rect -2966 57454 586890 57486
rect -2966 57218 -2934 57454
rect -2698 57218 -2614 57454
rect -2378 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 586302 57454
rect 586538 57218 586622 57454
rect 586858 57218 586890 57454
rect -2966 57134 586890 57218
rect -2966 56898 -2934 57134
rect -2698 56898 -2614 57134
rect -2378 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 586302 57134
rect 586538 56898 586622 57134
rect 586858 56898 586890 57134
rect -2966 56866 586890 56898
rect -8726 50614 592650 50646
rect -8726 50378 -7734 50614
rect -7498 50378 -7414 50614
rect -7178 50378 12986 50614
rect 13222 50378 13306 50614
rect 13542 50378 48986 50614
rect 49222 50378 49306 50614
rect 49542 50378 84986 50614
rect 85222 50378 85306 50614
rect 85542 50378 120986 50614
rect 121222 50378 121306 50614
rect 121542 50378 156986 50614
rect 157222 50378 157306 50614
rect 157542 50378 192986 50614
rect 193222 50378 193306 50614
rect 193542 50378 228986 50614
rect 229222 50378 229306 50614
rect 229542 50378 264986 50614
rect 265222 50378 265306 50614
rect 265542 50378 300986 50614
rect 301222 50378 301306 50614
rect 301542 50378 336986 50614
rect 337222 50378 337306 50614
rect 337542 50378 372986 50614
rect 373222 50378 373306 50614
rect 373542 50378 408986 50614
rect 409222 50378 409306 50614
rect 409542 50378 444986 50614
rect 445222 50378 445306 50614
rect 445542 50378 480986 50614
rect 481222 50378 481306 50614
rect 481542 50378 516986 50614
rect 517222 50378 517306 50614
rect 517542 50378 552986 50614
rect 553222 50378 553306 50614
rect 553542 50378 591102 50614
rect 591338 50378 591422 50614
rect 591658 50378 592650 50614
rect -8726 50294 592650 50378
rect -8726 50058 -7734 50294
rect -7498 50058 -7414 50294
rect -7178 50058 12986 50294
rect 13222 50058 13306 50294
rect 13542 50058 48986 50294
rect 49222 50058 49306 50294
rect 49542 50058 84986 50294
rect 85222 50058 85306 50294
rect 85542 50058 120986 50294
rect 121222 50058 121306 50294
rect 121542 50058 156986 50294
rect 157222 50058 157306 50294
rect 157542 50058 192986 50294
rect 193222 50058 193306 50294
rect 193542 50058 228986 50294
rect 229222 50058 229306 50294
rect 229542 50058 264986 50294
rect 265222 50058 265306 50294
rect 265542 50058 300986 50294
rect 301222 50058 301306 50294
rect 301542 50058 336986 50294
rect 337222 50058 337306 50294
rect 337542 50058 372986 50294
rect 373222 50058 373306 50294
rect 373542 50058 408986 50294
rect 409222 50058 409306 50294
rect 409542 50058 444986 50294
rect 445222 50058 445306 50294
rect 445542 50058 480986 50294
rect 481222 50058 481306 50294
rect 481542 50058 516986 50294
rect 517222 50058 517306 50294
rect 517542 50058 552986 50294
rect 553222 50058 553306 50294
rect 553542 50058 591102 50294
rect 591338 50058 591422 50294
rect 591658 50058 592650 50294
rect -8726 50026 592650 50058
rect -6806 46894 590730 46926
rect -6806 46658 -5814 46894
rect -5578 46658 -5494 46894
rect -5258 46658 9266 46894
rect 9502 46658 9586 46894
rect 9822 46658 45266 46894
rect 45502 46658 45586 46894
rect 45822 46658 81266 46894
rect 81502 46658 81586 46894
rect 81822 46658 117266 46894
rect 117502 46658 117586 46894
rect 117822 46658 153266 46894
rect 153502 46658 153586 46894
rect 153822 46658 189266 46894
rect 189502 46658 189586 46894
rect 189822 46658 225266 46894
rect 225502 46658 225586 46894
rect 225822 46658 261266 46894
rect 261502 46658 261586 46894
rect 261822 46658 297266 46894
rect 297502 46658 297586 46894
rect 297822 46658 333266 46894
rect 333502 46658 333586 46894
rect 333822 46658 369266 46894
rect 369502 46658 369586 46894
rect 369822 46658 405266 46894
rect 405502 46658 405586 46894
rect 405822 46658 441266 46894
rect 441502 46658 441586 46894
rect 441822 46658 477266 46894
rect 477502 46658 477586 46894
rect 477822 46658 513266 46894
rect 513502 46658 513586 46894
rect 513822 46658 549266 46894
rect 549502 46658 549586 46894
rect 549822 46658 589182 46894
rect 589418 46658 589502 46894
rect 589738 46658 590730 46894
rect -6806 46574 590730 46658
rect -6806 46338 -5814 46574
rect -5578 46338 -5494 46574
rect -5258 46338 9266 46574
rect 9502 46338 9586 46574
rect 9822 46338 45266 46574
rect 45502 46338 45586 46574
rect 45822 46338 81266 46574
rect 81502 46338 81586 46574
rect 81822 46338 117266 46574
rect 117502 46338 117586 46574
rect 117822 46338 153266 46574
rect 153502 46338 153586 46574
rect 153822 46338 189266 46574
rect 189502 46338 189586 46574
rect 189822 46338 225266 46574
rect 225502 46338 225586 46574
rect 225822 46338 261266 46574
rect 261502 46338 261586 46574
rect 261822 46338 297266 46574
rect 297502 46338 297586 46574
rect 297822 46338 333266 46574
rect 333502 46338 333586 46574
rect 333822 46338 369266 46574
rect 369502 46338 369586 46574
rect 369822 46338 405266 46574
rect 405502 46338 405586 46574
rect 405822 46338 441266 46574
rect 441502 46338 441586 46574
rect 441822 46338 477266 46574
rect 477502 46338 477586 46574
rect 477822 46338 513266 46574
rect 513502 46338 513586 46574
rect 513822 46338 549266 46574
rect 549502 46338 549586 46574
rect 549822 46338 589182 46574
rect 589418 46338 589502 46574
rect 589738 46338 590730 46574
rect -6806 46306 590730 46338
rect -4886 43174 588810 43206
rect -4886 42938 -3894 43174
rect -3658 42938 -3574 43174
rect -3338 42938 5546 43174
rect 5782 42938 5866 43174
rect 6102 42938 41546 43174
rect 41782 42938 41866 43174
rect 42102 42938 77546 43174
rect 77782 42938 77866 43174
rect 78102 42938 113546 43174
rect 113782 42938 113866 43174
rect 114102 42938 149546 43174
rect 149782 42938 149866 43174
rect 150102 42938 185546 43174
rect 185782 42938 185866 43174
rect 186102 42938 221546 43174
rect 221782 42938 221866 43174
rect 222102 42938 257546 43174
rect 257782 42938 257866 43174
rect 258102 42938 293546 43174
rect 293782 42938 293866 43174
rect 294102 42938 329546 43174
rect 329782 42938 329866 43174
rect 330102 42938 365546 43174
rect 365782 42938 365866 43174
rect 366102 42938 401546 43174
rect 401782 42938 401866 43174
rect 402102 42938 437546 43174
rect 437782 42938 437866 43174
rect 438102 42938 473546 43174
rect 473782 42938 473866 43174
rect 474102 42938 509546 43174
rect 509782 42938 509866 43174
rect 510102 42938 545546 43174
rect 545782 42938 545866 43174
rect 546102 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 587262 43174
rect 587498 42938 587582 43174
rect 587818 42938 588810 43174
rect -4886 42854 588810 42938
rect -4886 42618 -3894 42854
rect -3658 42618 -3574 42854
rect -3338 42618 5546 42854
rect 5782 42618 5866 42854
rect 6102 42618 41546 42854
rect 41782 42618 41866 42854
rect 42102 42618 77546 42854
rect 77782 42618 77866 42854
rect 78102 42618 113546 42854
rect 113782 42618 113866 42854
rect 114102 42618 149546 42854
rect 149782 42618 149866 42854
rect 150102 42618 185546 42854
rect 185782 42618 185866 42854
rect 186102 42618 221546 42854
rect 221782 42618 221866 42854
rect 222102 42618 257546 42854
rect 257782 42618 257866 42854
rect 258102 42618 293546 42854
rect 293782 42618 293866 42854
rect 294102 42618 329546 42854
rect 329782 42618 329866 42854
rect 330102 42618 365546 42854
rect 365782 42618 365866 42854
rect 366102 42618 401546 42854
rect 401782 42618 401866 42854
rect 402102 42618 437546 42854
rect 437782 42618 437866 42854
rect 438102 42618 473546 42854
rect 473782 42618 473866 42854
rect 474102 42618 509546 42854
rect 509782 42618 509866 42854
rect 510102 42618 545546 42854
rect 545782 42618 545866 42854
rect 546102 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 587262 42854
rect 587498 42618 587582 42854
rect 587818 42618 588810 42854
rect -4886 42586 588810 42618
rect -2966 39454 586890 39486
rect -2966 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 586890 39454
rect -2966 39134 586890 39218
rect -2966 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 586890 39134
rect -2966 38866 586890 38898
rect -8726 32614 592650 32646
rect -8726 32378 -8694 32614
rect -8458 32378 -8374 32614
rect -8138 32378 30986 32614
rect 31222 32378 31306 32614
rect 31542 32378 66986 32614
rect 67222 32378 67306 32614
rect 67542 32378 102986 32614
rect 103222 32378 103306 32614
rect 103542 32378 138986 32614
rect 139222 32378 139306 32614
rect 139542 32378 174986 32614
rect 175222 32378 175306 32614
rect 175542 32378 210986 32614
rect 211222 32378 211306 32614
rect 211542 32378 246986 32614
rect 247222 32378 247306 32614
rect 247542 32378 282986 32614
rect 283222 32378 283306 32614
rect 283542 32378 318986 32614
rect 319222 32378 319306 32614
rect 319542 32378 354986 32614
rect 355222 32378 355306 32614
rect 355542 32378 390986 32614
rect 391222 32378 391306 32614
rect 391542 32378 426986 32614
rect 427222 32378 427306 32614
rect 427542 32378 462986 32614
rect 463222 32378 463306 32614
rect 463542 32378 498986 32614
rect 499222 32378 499306 32614
rect 499542 32378 534986 32614
rect 535222 32378 535306 32614
rect 535542 32378 570986 32614
rect 571222 32378 571306 32614
rect 571542 32378 592062 32614
rect 592298 32378 592382 32614
rect 592618 32378 592650 32614
rect -8726 32294 592650 32378
rect -8726 32058 -8694 32294
rect -8458 32058 -8374 32294
rect -8138 32058 30986 32294
rect 31222 32058 31306 32294
rect 31542 32058 66986 32294
rect 67222 32058 67306 32294
rect 67542 32058 102986 32294
rect 103222 32058 103306 32294
rect 103542 32058 138986 32294
rect 139222 32058 139306 32294
rect 139542 32058 174986 32294
rect 175222 32058 175306 32294
rect 175542 32058 210986 32294
rect 211222 32058 211306 32294
rect 211542 32058 246986 32294
rect 247222 32058 247306 32294
rect 247542 32058 282986 32294
rect 283222 32058 283306 32294
rect 283542 32058 318986 32294
rect 319222 32058 319306 32294
rect 319542 32058 354986 32294
rect 355222 32058 355306 32294
rect 355542 32058 390986 32294
rect 391222 32058 391306 32294
rect 391542 32058 426986 32294
rect 427222 32058 427306 32294
rect 427542 32058 462986 32294
rect 463222 32058 463306 32294
rect 463542 32058 498986 32294
rect 499222 32058 499306 32294
rect 499542 32058 534986 32294
rect 535222 32058 535306 32294
rect 535542 32058 570986 32294
rect 571222 32058 571306 32294
rect 571542 32058 592062 32294
rect 592298 32058 592382 32294
rect 592618 32058 592650 32294
rect -8726 32026 592650 32058
rect -6806 28894 590730 28926
rect -6806 28658 -6774 28894
rect -6538 28658 -6454 28894
rect -6218 28658 27266 28894
rect 27502 28658 27586 28894
rect 27822 28658 63266 28894
rect 63502 28658 63586 28894
rect 63822 28658 99266 28894
rect 99502 28658 99586 28894
rect 99822 28658 135266 28894
rect 135502 28658 135586 28894
rect 135822 28658 171266 28894
rect 171502 28658 171586 28894
rect 171822 28658 207266 28894
rect 207502 28658 207586 28894
rect 207822 28658 243266 28894
rect 243502 28658 243586 28894
rect 243822 28658 279266 28894
rect 279502 28658 279586 28894
rect 279822 28658 315266 28894
rect 315502 28658 315586 28894
rect 315822 28658 351266 28894
rect 351502 28658 351586 28894
rect 351822 28658 387266 28894
rect 387502 28658 387586 28894
rect 387822 28658 423266 28894
rect 423502 28658 423586 28894
rect 423822 28658 459266 28894
rect 459502 28658 459586 28894
rect 459822 28658 495266 28894
rect 495502 28658 495586 28894
rect 495822 28658 531266 28894
rect 531502 28658 531586 28894
rect 531822 28658 567266 28894
rect 567502 28658 567586 28894
rect 567822 28658 590142 28894
rect 590378 28658 590462 28894
rect 590698 28658 590730 28894
rect -6806 28574 590730 28658
rect -6806 28338 -6774 28574
rect -6538 28338 -6454 28574
rect -6218 28338 27266 28574
rect 27502 28338 27586 28574
rect 27822 28338 63266 28574
rect 63502 28338 63586 28574
rect 63822 28338 99266 28574
rect 99502 28338 99586 28574
rect 99822 28338 135266 28574
rect 135502 28338 135586 28574
rect 135822 28338 171266 28574
rect 171502 28338 171586 28574
rect 171822 28338 207266 28574
rect 207502 28338 207586 28574
rect 207822 28338 243266 28574
rect 243502 28338 243586 28574
rect 243822 28338 279266 28574
rect 279502 28338 279586 28574
rect 279822 28338 315266 28574
rect 315502 28338 315586 28574
rect 315822 28338 351266 28574
rect 351502 28338 351586 28574
rect 351822 28338 387266 28574
rect 387502 28338 387586 28574
rect 387822 28338 423266 28574
rect 423502 28338 423586 28574
rect 423822 28338 459266 28574
rect 459502 28338 459586 28574
rect 459822 28338 495266 28574
rect 495502 28338 495586 28574
rect 495822 28338 531266 28574
rect 531502 28338 531586 28574
rect 531822 28338 567266 28574
rect 567502 28338 567586 28574
rect 567822 28338 590142 28574
rect 590378 28338 590462 28574
rect 590698 28338 590730 28574
rect -6806 28306 590730 28338
rect -4886 25174 588810 25206
rect -4886 24938 -4854 25174
rect -4618 24938 -4534 25174
rect -4298 24938 23546 25174
rect 23782 24938 23866 25174
rect 24102 24938 59546 25174
rect 59782 24938 59866 25174
rect 60102 24938 95546 25174
rect 95782 24938 95866 25174
rect 96102 24938 131546 25174
rect 131782 24938 131866 25174
rect 132102 24938 167546 25174
rect 167782 24938 167866 25174
rect 168102 24938 203546 25174
rect 203782 24938 203866 25174
rect 204102 24938 239546 25174
rect 239782 24938 239866 25174
rect 240102 24938 275546 25174
rect 275782 24938 275866 25174
rect 276102 24938 311546 25174
rect 311782 24938 311866 25174
rect 312102 24938 347546 25174
rect 347782 24938 347866 25174
rect 348102 24938 383546 25174
rect 383782 24938 383866 25174
rect 384102 24938 419546 25174
rect 419782 24938 419866 25174
rect 420102 24938 455546 25174
rect 455782 24938 455866 25174
rect 456102 24938 491546 25174
rect 491782 24938 491866 25174
rect 492102 24938 527546 25174
rect 527782 24938 527866 25174
rect 528102 24938 563546 25174
rect 563782 24938 563866 25174
rect 564102 24938 588222 25174
rect 588458 24938 588542 25174
rect 588778 24938 588810 25174
rect -4886 24854 588810 24938
rect -4886 24618 -4854 24854
rect -4618 24618 -4534 24854
rect -4298 24618 23546 24854
rect 23782 24618 23866 24854
rect 24102 24618 59546 24854
rect 59782 24618 59866 24854
rect 60102 24618 95546 24854
rect 95782 24618 95866 24854
rect 96102 24618 131546 24854
rect 131782 24618 131866 24854
rect 132102 24618 167546 24854
rect 167782 24618 167866 24854
rect 168102 24618 203546 24854
rect 203782 24618 203866 24854
rect 204102 24618 239546 24854
rect 239782 24618 239866 24854
rect 240102 24618 275546 24854
rect 275782 24618 275866 24854
rect 276102 24618 311546 24854
rect 311782 24618 311866 24854
rect 312102 24618 347546 24854
rect 347782 24618 347866 24854
rect 348102 24618 383546 24854
rect 383782 24618 383866 24854
rect 384102 24618 419546 24854
rect 419782 24618 419866 24854
rect 420102 24618 455546 24854
rect 455782 24618 455866 24854
rect 456102 24618 491546 24854
rect 491782 24618 491866 24854
rect 492102 24618 527546 24854
rect 527782 24618 527866 24854
rect 528102 24618 563546 24854
rect 563782 24618 563866 24854
rect 564102 24618 588222 24854
rect 588458 24618 588542 24854
rect 588778 24618 588810 24854
rect -4886 24586 588810 24618
rect -2966 21454 586890 21486
rect -2966 21218 -2934 21454
rect -2698 21218 -2614 21454
rect -2378 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 586302 21454
rect 586538 21218 586622 21454
rect 586858 21218 586890 21454
rect -2966 21134 586890 21218
rect -2966 20898 -2934 21134
rect -2698 20898 -2614 21134
rect -2378 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 586302 21134
rect 586538 20898 586622 21134
rect 586858 20898 586890 21134
rect -2966 20866 586890 20898
rect -8726 14614 592650 14646
rect -8726 14378 -7734 14614
rect -7498 14378 -7414 14614
rect -7178 14378 12986 14614
rect 13222 14378 13306 14614
rect 13542 14378 48986 14614
rect 49222 14378 49306 14614
rect 49542 14378 84986 14614
rect 85222 14378 85306 14614
rect 85542 14378 120986 14614
rect 121222 14378 121306 14614
rect 121542 14378 156986 14614
rect 157222 14378 157306 14614
rect 157542 14378 192986 14614
rect 193222 14378 193306 14614
rect 193542 14378 228986 14614
rect 229222 14378 229306 14614
rect 229542 14378 264986 14614
rect 265222 14378 265306 14614
rect 265542 14378 300986 14614
rect 301222 14378 301306 14614
rect 301542 14378 336986 14614
rect 337222 14378 337306 14614
rect 337542 14378 372986 14614
rect 373222 14378 373306 14614
rect 373542 14378 408986 14614
rect 409222 14378 409306 14614
rect 409542 14378 444986 14614
rect 445222 14378 445306 14614
rect 445542 14378 480986 14614
rect 481222 14378 481306 14614
rect 481542 14378 516986 14614
rect 517222 14378 517306 14614
rect 517542 14378 552986 14614
rect 553222 14378 553306 14614
rect 553542 14378 591102 14614
rect 591338 14378 591422 14614
rect 591658 14378 592650 14614
rect -8726 14294 592650 14378
rect -8726 14058 -7734 14294
rect -7498 14058 -7414 14294
rect -7178 14058 12986 14294
rect 13222 14058 13306 14294
rect 13542 14058 48986 14294
rect 49222 14058 49306 14294
rect 49542 14058 84986 14294
rect 85222 14058 85306 14294
rect 85542 14058 120986 14294
rect 121222 14058 121306 14294
rect 121542 14058 156986 14294
rect 157222 14058 157306 14294
rect 157542 14058 192986 14294
rect 193222 14058 193306 14294
rect 193542 14058 228986 14294
rect 229222 14058 229306 14294
rect 229542 14058 264986 14294
rect 265222 14058 265306 14294
rect 265542 14058 300986 14294
rect 301222 14058 301306 14294
rect 301542 14058 336986 14294
rect 337222 14058 337306 14294
rect 337542 14058 372986 14294
rect 373222 14058 373306 14294
rect 373542 14058 408986 14294
rect 409222 14058 409306 14294
rect 409542 14058 444986 14294
rect 445222 14058 445306 14294
rect 445542 14058 480986 14294
rect 481222 14058 481306 14294
rect 481542 14058 516986 14294
rect 517222 14058 517306 14294
rect 517542 14058 552986 14294
rect 553222 14058 553306 14294
rect 553542 14058 591102 14294
rect 591338 14058 591422 14294
rect 591658 14058 592650 14294
rect -8726 14026 592650 14058
rect -6806 10894 590730 10926
rect -6806 10658 -5814 10894
rect -5578 10658 -5494 10894
rect -5258 10658 9266 10894
rect 9502 10658 9586 10894
rect 9822 10658 45266 10894
rect 45502 10658 45586 10894
rect 45822 10658 81266 10894
rect 81502 10658 81586 10894
rect 81822 10658 117266 10894
rect 117502 10658 117586 10894
rect 117822 10658 153266 10894
rect 153502 10658 153586 10894
rect 153822 10658 189266 10894
rect 189502 10658 189586 10894
rect 189822 10658 225266 10894
rect 225502 10658 225586 10894
rect 225822 10658 261266 10894
rect 261502 10658 261586 10894
rect 261822 10658 297266 10894
rect 297502 10658 297586 10894
rect 297822 10658 333266 10894
rect 333502 10658 333586 10894
rect 333822 10658 369266 10894
rect 369502 10658 369586 10894
rect 369822 10658 405266 10894
rect 405502 10658 405586 10894
rect 405822 10658 441266 10894
rect 441502 10658 441586 10894
rect 441822 10658 477266 10894
rect 477502 10658 477586 10894
rect 477822 10658 513266 10894
rect 513502 10658 513586 10894
rect 513822 10658 549266 10894
rect 549502 10658 549586 10894
rect 549822 10658 589182 10894
rect 589418 10658 589502 10894
rect 589738 10658 590730 10894
rect -6806 10574 590730 10658
rect -6806 10338 -5814 10574
rect -5578 10338 -5494 10574
rect -5258 10338 9266 10574
rect 9502 10338 9586 10574
rect 9822 10338 45266 10574
rect 45502 10338 45586 10574
rect 45822 10338 81266 10574
rect 81502 10338 81586 10574
rect 81822 10338 117266 10574
rect 117502 10338 117586 10574
rect 117822 10338 153266 10574
rect 153502 10338 153586 10574
rect 153822 10338 189266 10574
rect 189502 10338 189586 10574
rect 189822 10338 225266 10574
rect 225502 10338 225586 10574
rect 225822 10338 261266 10574
rect 261502 10338 261586 10574
rect 261822 10338 297266 10574
rect 297502 10338 297586 10574
rect 297822 10338 333266 10574
rect 333502 10338 333586 10574
rect 333822 10338 369266 10574
rect 369502 10338 369586 10574
rect 369822 10338 405266 10574
rect 405502 10338 405586 10574
rect 405822 10338 441266 10574
rect 441502 10338 441586 10574
rect 441822 10338 477266 10574
rect 477502 10338 477586 10574
rect 477822 10338 513266 10574
rect 513502 10338 513586 10574
rect 513822 10338 549266 10574
rect 549502 10338 549586 10574
rect 549822 10338 589182 10574
rect 589418 10338 589502 10574
rect 589738 10338 590730 10574
rect -6806 10306 590730 10338
rect -4886 7174 588810 7206
rect -4886 6938 -3894 7174
rect -3658 6938 -3574 7174
rect -3338 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 41546 7174
rect 41782 6938 41866 7174
rect 42102 6938 77546 7174
rect 77782 6938 77866 7174
rect 78102 6938 113546 7174
rect 113782 6938 113866 7174
rect 114102 6938 149546 7174
rect 149782 6938 149866 7174
rect 150102 6938 185546 7174
rect 185782 6938 185866 7174
rect 186102 6938 221546 7174
rect 221782 6938 221866 7174
rect 222102 6938 257546 7174
rect 257782 6938 257866 7174
rect 258102 6938 293546 7174
rect 293782 6938 293866 7174
rect 294102 6938 329546 7174
rect 329782 6938 329866 7174
rect 330102 6938 365546 7174
rect 365782 6938 365866 7174
rect 366102 6938 401546 7174
rect 401782 6938 401866 7174
rect 402102 6938 437546 7174
rect 437782 6938 437866 7174
rect 438102 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 509546 7174
rect 509782 6938 509866 7174
rect 510102 6938 545546 7174
rect 545782 6938 545866 7174
rect 546102 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 587262 7174
rect 587498 6938 587582 7174
rect 587818 6938 588810 7174
rect -4886 6854 588810 6938
rect -4886 6618 -3894 6854
rect -3658 6618 -3574 6854
rect -3338 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 41546 6854
rect 41782 6618 41866 6854
rect 42102 6618 77546 6854
rect 77782 6618 77866 6854
rect 78102 6618 113546 6854
rect 113782 6618 113866 6854
rect 114102 6618 149546 6854
rect 149782 6618 149866 6854
rect 150102 6618 185546 6854
rect 185782 6618 185866 6854
rect 186102 6618 221546 6854
rect 221782 6618 221866 6854
rect 222102 6618 257546 6854
rect 257782 6618 257866 6854
rect 258102 6618 293546 6854
rect 293782 6618 293866 6854
rect 294102 6618 329546 6854
rect 329782 6618 329866 6854
rect 330102 6618 365546 6854
rect 365782 6618 365866 6854
rect 366102 6618 401546 6854
rect 401782 6618 401866 6854
rect 402102 6618 437546 6854
rect 437782 6618 437866 6854
rect 438102 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 509546 6854
rect 509782 6618 509866 6854
rect 510102 6618 545546 6854
rect 545782 6618 545866 6854
rect 546102 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 587262 6854
rect 587498 6618 587582 6854
rect 587818 6618 588810 6854
rect -4886 6586 588810 6618
rect -2966 3454 586890 3486
rect -2966 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 586890 3454
rect -2966 3134 586890 3218
rect -2966 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 586890 3134
rect -2966 2866 586890 2898
rect -2006 -346 585930 -314
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect -2006 -666 585930 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect -2006 -934 585930 -902
rect -2966 -1306 586890 -1274
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 19826 -1306
rect 20062 -1542 20146 -1306
rect 20382 -1542 55826 -1306
rect 56062 -1542 56146 -1306
rect 56382 -1542 91826 -1306
rect 92062 -1542 92146 -1306
rect 92382 -1542 127826 -1306
rect 128062 -1542 128146 -1306
rect 128382 -1542 163826 -1306
rect 164062 -1542 164146 -1306
rect 164382 -1542 199826 -1306
rect 200062 -1542 200146 -1306
rect 200382 -1542 235826 -1306
rect 236062 -1542 236146 -1306
rect 236382 -1542 271826 -1306
rect 272062 -1542 272146 -1306
rect 272382 -1542 307826 -1306
rect 308062 -1542 308146 -1306
rect 308382 -1542 343826 -1306
rect 344062 -1542 344146 -1306
rect 344382 -1542 379826 -1306
rect 380062 -1542 380146 -1306
rect 380382 -1542 415826 -1306
rect 416062 -1542 416146 -1306
rect 416382 -1542 451826 -1306
rect 452062 -1542 452146 -1306
rect 452382 -1542 487826 -1306
rect 488062 -1542 488146 -1306
rect 488382 -1542 523826 -1306
rect 524062 -1542 524146 -1306
rect 524382 -1542 559826 -1306
rect 560062 -1542 560146 -1306
rect 560382 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect -2966 -1626 586890 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 19826 -1626
rect 20062 -1862 20146 -1626
rect 20382 -1862 55826 -1626
rect 56062 -1862 56146 -1626
rect 56382 -1862 91826 -1626
rect 92062 -1862 92146 -1626
rect 92382 -1862 127826 -1626
rect 128062 -1862 128146 -1626
rect 128382 -1862 163826 -1626
rect 164062 -1862 164146 -1626
rect 164382 -1862 199826 -1626
rect 200062 -1862 200146 -1626
rect 200382 -1862 235826 -1626
rect 236062 -1862 236146 -1626
rect 236382 -1862 271826 -1626
rect 272062 -1862 272146 -1626
rect 272382 -1862 307826 -1626
rect 308062 -1862 308146 -1626
rect 308382 -1862 343826 -1626
rect 344062 -1862 344146 -1626
rect 344382 -1862 379826 -1626
rect 380062 -1862 380146 -1626
rect 380382 -1862 415826 -1626
rect 416062 -1862 416146 -1626
rect 416382 -1862 451826 -1626
rect 452062 -1862 452146 -1626
rect 452382 -1862 487826 -1626
rect 488062 -1862 488146 -1626
rect 488382 -1862 523826 -1626
rect 524062 -1862 524146 -1626
rect 524382 -1862 559826 -1626
rect 560062 -1862 560146 -1626
rect 560382 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect -2966 -1894 586890 -1862
rect -3926 -2266 587850 -2234
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 5546 -2266
rect 5782 -2502 5866 -2266
rect 6102 -2502 41546 -2266
rect 41782 -2502 41866 -2266
rect 42102 -2502 77546 -2266
rect 77782 -2502 77866 -2266
rect 78102 -2502 113546 -2266
rect 113782 -2502 113866 -2266
rect 114102 -2502 149546 -2266
rect 149782 -2502 149866 -2266
rect 150102 -2502 185546 -2266
rect 185782 -2502 185866 -2266
rect 186102 -2502 221546 -2266
rect 221782 -2502 221866 -2266
rect 222102 -2502 257546 -2266
rect 257782 -2502 257866 -2266
rect 258102 -2502 293546 -2266
rect 293782 -2502 293866 -2266
rect 294102 -2502 329546 -2266
rect 329782 -2502 329866 -2266
rect 330102 -2502 365546 -2266
rect 365782 -2502 365866 -2266
rect 366102 -2502 401546 -2266
rect 401782 -2502 401866 -2266
rect 402102 -2502 437546 -2266
rect 437782 -2502 437866 -2266
rect 438102 -2502 473546 -2266
rect 473782 -2502 473866 -2266
rect 474102 -2502 509546 -2266
rect 509782 -2502 509866 -2266
rect 510102 -2502 545546 -2266
rect 545782 -2502 545866 -2266
rect 546102 -2502 581546 -2266
rect 581782 -2502 581866 -2266
rect 582102 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect -3926 -2586 587850 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 5546 -2586
rect 5782 -2822 5866 -2586
rect 6102 -2822 41546 -2586
rect 41782 -2822 41866 -2586
rect 42102 -2822 77546 -2586
rect 77782 -2822 77866 -2586
rect 78102 -2822 113546 -2586
rect 113782 -2822 113866 -2586
rect 114102 -2822 149546 -2586
rect 149782 -2822 149866 -2586
rect 150102 -2822 185546 -2586
rect 185782 -2822 185866 -2586
rect 186102 -2822 221546 -2586
rect 221782 -2822 221866 -2586
rect 222102 -2822 257546 -2586
rect 257782 -2822 257866 -2586
rect 258102 -2822 293546 -2586
rect 293782 -2822 293866 -2586
rect 294102 -2822 329546 -2586
rect 329782 -2822 329866 -2586
rect 330102 -2822 365546 -2586
rect 365782 -2822 365866 -2586
rect 366102 -2822 401546 -2586
rect 401782 -2822 401866 -2586
rect 402102 -2822 437546 -2586
rect 437782 -2822 437866 -2586
rect 438102 -2822 473546 -2586
rect 473782 -2822 473866 -2586
rect 474102 -2822 509546 -2586
rect 509782 -2822 509866 -2586
rect 510102 -2822 545546 -2586
rect 545782 -2822 545866 -2586
rect 546102 -2822 581546 -2586
rect 581782 -2822 581866 -2586
rect 582102 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect -3926 -2854 587850 -2822
rect -4886 -3226 588810 -3194
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 23546 -3226
rect 23782 -3462 23866 -3226
rect 24102 -3462 59546 -3226
rect 59782 -3462 59866 -3226
rect 60102 -3462 95546 -3226
rect 95782 -3462 95866 -3226
rect 96102 -3462 131546 -3226
rect 131782 -3462 131866 -3226
rect 132102 -3462 167546 -3226
rect 167782 -3462 167866 -3226
rect 168102 -3462 203546 -3226
rect 203782 -3462 203866 -3226
rect 204102 -3462 239546 -3226
rect 239782 -3462 239866 -3226
rect 240102 -3462 275546 -3226
rect 275782 -3462 275866 -3226
rect 276102 -3462 311546 -3226
rect 311782 -3462 311866 -3226
rect 312102 -3462 347546 -3226
rect 347782 -3462 347866 -3226
rect 348102 -3462 383546 -3226
rect 383782 -3462 383866 -3226
rect 384102 -3462 419546 -3226
rect 419782 -3462 419866 -3226
rect 420102 -3462 455546 -3226
rect 455782 -3462 455866 -3226
rect 456102 -3462 491546 -3226
rect 491782 -3462 491866 -3226
rect 492102 -3462 527546 -3226
rect 527782 -3462 527866 -3226
rect 528102 -3462 563546 -3226
rect 563782 -3462 563866 -3226
rect 564102 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect -4886 -3546 588810 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 23546 -3546
rect 23782 -3782 23866 -3546
rect 24102 -3782 59546 -3546
rect 59782 -3782 59866 -3546
rect 60102 -3782 95546 -3546
rect 95782 -3782 95866 -3546
rect 96102 -3782 131546 -3546
rect 131782 -3782 131866 -3546
rect 132102 -3782 167546 -3546
rect 167782 -3782 167866 -3546
rect 168102 -3782 203546 -3546
rect 203782 -3782 203866 -3546
rect 204102 -3782 239546 -3546
rect 239782 -3782 239866 -3546
rect 240102 -3782 275546 -3546
rect 275782 -3782 275866 -3546
rect 276102 -3782 311546 -3546
rect 311782 -3782 311866 -3546
rect 312102 -3782 347546 -3546
rect 347782 -3782 347866 -3546
rect 348102 -3782 383546 -3546
rect 383782 -3782 383866 -3546
rect 384102 -3782 419546 -3546
rect 419782 -3782 419866 -3546
rect 420102 -3782 455546 -3546
rect 455782 -3782 455866 -3546
rect 456102 -3782 491546 -3546
rect 491782 -3782 491866 -3546
rect 492102 -3782 527546 -3546
rect 527782 -3782 527866 -3546
rect 528102 -3782 563546 -3546
rect 563782 -3782 563866 -3546
rect 564102 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect -4886 -3814 588810 -3782
rect -5846 -4186 589770 -4154
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 9266 -4186
rect 9502 -4422 9586 -4186
rect 9822 -4422 45266 -4186
rect 45502 -4422 45586 -4186
rect 45822 -4422 81266 -4186
rect 81502 -4422 81586 -4186
rect 81822 -4422 117266 -4186
rect 117502 -4422 117586 -4186
rect 117822 -4422 153266 -4186
rect 153502 -4422 153586 -4186
rect 153822 -4422 189266 -4186
rect 189502 -4422 189586 -4186
rect 189822 -4422 225266 -4186
rect 225502 -4422 225586 -4186
rect 225822 -4422 261266 -4186
rect 261502 -4422 261586 -4186
rect 261822 -4422 297266 -4186
rect 297502 -4422 297586 -4186
rect 297822 -4422 333266 -4186
rect 333502 -4422 333586 -4186
rect 333822 -4422 369266 -4186
rect 369502 -4422 369586 -4186
rect 369822 -4422 405266 -4186
rect 405502 -4422 405586 -4186
rect 405822 -4422 441266 -4186
rect 441502 -4422 441586 -4186
rect 441822 -4422 477266 -4186
rect 477502 -4422 477586 -4186
rect 477822 -4422 513266 -4186
rect 513502 -4422 513586 -4186
rect 513822 -4422 549266 -4186
rect 549502 -4422 549586 -4186
rect 549822 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect -5846 -4506 589770 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 9266 -4506
rect 9502 -4742 9586 -4506
rect 9822 -4742 45266 -4506
rect 45502 -4742 45586 -4506
rect 45822 -4742 81266 -4506
rect 81502 -4742 81586 -4506
rect 81822 -4742 117266 -4506
rect 117502 -4742 117586 -4506
rect 117822 -4742 153266 -4506
rect 153502 -4742 153586 -4506
rect 153822 -4742 189266 -4506
rect 189502 -4742 189586 -4506
rect 189822 -4742 225266 -4506
rect 225502 -4742 225586 -4506
rect 225822 -4742 261266 -4506
rect 261502 -4742 261586 -4506
rect 261822 -4742 297266 -4506
rect 297502 -4742 297586 -4506
rect 297822 -4742 333266 -4506
rect 333502 -4742 333586 -4506
rect 333822 -4742 369266 -4506
rect 369502 -4742 369586 -4506
rect 369822 -4742 405266 -4506
rect 405502 -4742 405586 -4506
rect 405822 -4742 441266 -4506
rect 441502 -4742 441586 -4506
rect 441822 -4742 477266 -4506
rect 477502 -4742 477586 -4506
rect 477822 -4742 513266 -4506
rect 513502 -4742 513586 -4506
rect 513822 -4742 549266 -4506
rect 549502 -4742 549586 -4506
rect 549822 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect -5846 -4774 589770 -4742
rect -6806 -5146 590730 -5114
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 27266 -5146
rect 27502 -5382 27586 -5146
rect 27822 -5382 63266 -5146
rect 63502 -5382 63586 -5146
rect 63822 -5382 99266 -5146
rect 99502 -5382 99586 -5146
rect 99822 -5382 135266 -5146
rect 135502 -5382 135586 -5146
rect 135822 -5382 171266 -5146
rect 171502 -5382 171586 -5146
rect 171822 -5382 207266 -5146
rect 207502 -5382 207586 -5146
rect 207822 -5382 243266 -5146
rect 243502 -5382 243586 -5146
rect 243822 -5382 279266 -5146
rect 279502 -5382 279586 -5146
rect 279822 -5382 315266 -5146
rect 315502 -5382 315586 -5146
rect 315822 -5382 351266 -5146
rect 351502 -5382 351586 -5146
rect 351822 -5382 387266 -5146
rect 387502 -5382 387586 -5146
rect 387822 -5382 423266 -5146
rect 423502 -5382 423586 -5146
rect 423822 -5382 459266 -5146
rect 459502 -5382 459586 -5146
rect 459822 -5382 495266 -5146
rect 495502 -5382 495586 -5146
rect 495822 -5382 531266 -5146
rect 531502 -5382 531586 -5146
rect 531822 -5382 567266 -5146
rect 567502 -5382 567586 -5146
rect 567822 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect -6806 -5466 590730 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 27266 -5466
rect 27502 -5702 27586 -5466
rect 27822 -5702 63266 -5466
rect 63502 -5702 63586 -5466
rect 63822 -5702 99266 -5466
rect 99502 -5702 99586 -5466
rect 99822 -5702 135266 -5466
rect 135502 -5702 135586 -5466
rect 135822 -5702 171266 -5466
rect 171502 -5702 171586 -5466
rect 171822 -5702 207266 -5466
rect 207502 -5702 207586 -5466
rect 207822 -5702 243266 -5466
rect 243502 -5702 243586 -5466
rect 243822 -5702 279266 -5466
rect 279502 -5702 279586 -5466
rect 279822 -5702 315266 -5466
rect 315502 -5702 315586 -5466
rect 315822 -5702 351266 -5466
rect 351502 -5702 351586 -5466
rect 351822 -5702 387266 -5466
rect 387502 -5702 387586 -5466
rect 387822 -5702 423266 -5466
rect 423502 -5702 423586 -5466
rect 423822 -5702 459266 -5466
rect 459502 -5702 459586 -5466
rect 459822 -5702 495266 -5466
rect 495502 -5702 495586 -5466
rect 495822 -5702 531266 -5466
rect 531502 -5702 531586 -5466
rect 531822 -5702 567266 -5466
rect 567502 -5702 567586 -5466
rect 567822 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect -6806 -5734 590730 -5702
rect -7766 -6106 591690 -6074
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 12986 -6106
rect 13222 -6342 13306 -6106
rect 13542 -6342 48986 -6106
rect 49222 -6342 49306 -6106
rect 49542 -6342 84986 -6106
rect 85222 -6342 85306 -6106
rect 85542 -6342 120986 -6106
rect 121222 -6342 121306 -6106
rect 121542 -6342 156986 -6106
rect 157222 -6342 157306 -6106
rect 157542 -6342 192986 -6106
rect 193222 -6342 193306 -6106
rect 193542 -6342 228986 -6106
rect 229222 -6342 229306 -6106
rect 229542 -6342 264986 -6106
rect 265222 -6342 265306 -6106
rect 265542 -6342 300986 -6106
rect 301222 -6342 301306 -6106
rect 301542 -6342 336986 -6106
rect 337222 -6342 337306 -6106
rect 337542 -6342 372986 -6106
rect 373222 -6342 373306 -6106
rect 373542 -6342 408986 -6106
rect 409222 -6342 409306 -6106
rect 409542 -6342 444986 -6106
rect 445222 -6342 445306 -6106
rect 445542 -6342 480986 -6106
rect 481222 -6342 481306 -6106
rect 481542 -6342 516986 -6106
rect 517222 -6342 517306 -6106
rect 517542 -6342 552986 -6106
rect 553222 -6342 553306 -6106
rect 553542 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect -7766 -6426 591690 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 12986 -6426
rect 13222 -6662 13306 -6426
rect 13542 -6662 48986 -6426
rect 49222 -6662 49306 -6426
rect 49542 -6662 84986 -6426
rect 85222 -6662 85306 -6426
rect 85542 -6662 120986 -6426
rect 121222 -6662 121306 -6426
rect 121542 -6662 156986 -6426
rect 157222 -6662 157306 -6426
rect 157542 -6662 192986 -6426
rect 193222 -6662 193306 -6426
rect 193542 -6662 228986 -6426
rect 229222 -6662 229306 -6426
rect 229542 -6662 264986 -6426
rect 265222 -6662 265306 -6426
rect 265542 -6662 300986 -6426
rect 301222 -6662 301306 -6426
rect 301542 -6662 336986 -6426
rect 337222 -6662 337306 -6426
rect 337542 -6662 372986 -6426
rect 373222 -6662 373306 -6426
rect 373542 -6662 408986 -6426
rect 409222 -6662 409306 -6426
rect 409542 -6662 444986 -6426
rect 445222 -6662 445306 -6426
rect 445542 -6662 480986 -6426
rect 481222 -6662 481306 -6426
rect 481542 -6662 516986 -6426
rect 517222 -6662 517306 -6426
rect 517542 -6662 552986 -6426
rect 553222 -6662 553306 -6426
rect 553542 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect -7766 -6694 591690 -6662
rect -8726 -7066 592650 -7034
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 30986 -7066
rect 31222 -7302 31306 -7066
rect 31542 -7302 66986 -7066
rect 67222 -7302 67306 -7066
rect 67542 -7302 102986 -7066
rect 103222 -7302 103306 -7066
rect 103542 -7302 138986 -7066
rect 139222 -7302 139306 -7066
rect 139542 -7302 174986 -7066
rect 175222 -7302 175306 -7066
rect 175542 -7302 210986 -7066
rect 211222 -7302 211306 -7066
rect 211542 -7302 246986 -7066
rect 247222 -7302 247306 -7066
rect 247542 -7302 282986 -7066
rect 283222 -7302 283306 -7066
rect 283542 -7302 318986 -7066
rect 319222 -7302 319306 -7066
rect 319542 -7302 354986 -7066
rect 355222 -7302 355306 -7066
rect 355542 -7302 390986 -7066
rect 391222 -7302 391306 -7066
rect 391542 -7302 426986 -7066
rect 427222 -7302 427306 -7066
rect 427542 -7302 462986 -7066
rect 463222 -7302 463306 -7066
rect 463542 -7302 498986 -7066
rect 499222 -7302 499306 -7066
rect 499542 -7302 534986 -7066
rect 535222 -7302 535306 -7066
rect 535542 -7302 570986 -7066
rect 571222 -7302 571306 -7066
rect 571542 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect -8726 -7386 592650 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 30986 -7386
rect 31222 -7622 31306 -7386
rect 31542 -7622 66986 -7386
rect 67222 -7622 67306 -7386
rect 67542 -7622 102986 -7386
rect 103222 -7622 103306 -7386
rect 103542 -7622 138986 -7386
rect 139222 -7622 139306 -7386
rect 139542 -7622 174986 -7386
rect 175222 -7622 175306 -7386
rect 175542 -7622 210986 -7386
rect 211222 -7622 211306 -7386
rect 211542 -7622 246986 -7386
rect 247222 -7622 247306 -7386
rect 247542 -7622 282986 -7386
rect 283222 -7622 283306 -7386
rect 283542 -7622 318986 -7386
rect 319222 -7622 319306 -7386
rect 319542 -7622 354986 -7386
rect 355222 -7622 355306 -7386
rect 355542 -7622 390986 -7386
rect 391222 -7622 391306 -7386
rect 391542 -7622 426986 -7386
rect 427222 -7622 427306 -7386
rect 427542 -7622 462986 -7386
rect 463222 -7622 463306 -7386
rect 463542 -7622 498986 -7386
rect 499222 -7622 499306 -7386
rect 499542 -7622 534986 -7386
rect 535222 -7622 535306 -7386
rect 535542 -7622 570986 -7386
rect 571222 -7622 571306 -7386
rect 571542 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect -8726 -7654 592650 -7622
use user_project  mprj
timestamp 1647846298
transform 1 0 165800 0 1 200800
box 198 0 254274 307139
<< labels >>
rlabel metal3 s 583520 285276 584960 285516 6 analog_io[0]
port 0 nsew signal bidirectional
rlabel metal2 s 446098 703520 446210 704960 6 analog_io[10]
port 1 nsew signal bidirectional
rlabel metal2 s 381146 703520 381258 704960 6 analog_io[11]
port 2 nsew signal bidirectional
rlabel metal2 s 316286 703520 316398 704960 6 analog_io[12]
port 3 nsew signal bidirectional
rlabel metal2 s 251426 703520 251538 704960 6 analog_io[13]
port 4 nsew signal bidirectional
rlabel metal2 s 186474 703520 186586 704960 6 analog_io[14]
port 5 nsew signal bidirectional
rlabel metal2 s 121614 703520 121726 704960 6 analog_io[15]
port 6 nsew signal bidirectional
rlabel metal2 s 56754 703520 56866 704960 6 analog_io[16]
port 7 nsew signal bidirectional
rlabel metal3 s -960 697220 480 697460 4 analog_io[17]
port 8 nsew signal bidirectional
rlabel metal3 s -960 644996 480 645236 4 analog_io[18]
port 9 nsew signal bidirectional
rlabel metal3 s -960 592908 480 593148 4 analog_io[19]
port 10 nsew signal bidirectional
rlabel metal3 s 583520 338452 584960 338692 6 analog_io[1]
port 11 nsew signal bidirectional
rlabel metal3 s -960 540684 480 540924 4 analog_io[20]
port 12 nsew signal bidirectional
rlabel metal3 s -960 488596 480 488836 4 analog_io[21]
port 13 nsew signal bidirectional
rlabel metal3 s -960 436508 480 436748 4 analog_io[22]
port 14 nsew signal bidirectional
rlabel metal3 s -960 384284 480 384524 4 analog_io[23]
port 15 nsew signal bidirectional
rlabel metal3 s -960 332196 480 332436 4 analog_io[24]
port 16 nsew signal bidirectional
rlabel metal3 s -960 279972 480 280212 4 analog_io[25]
port 17 nsew signal bidirectional
rlabel metal3 s -960 227884 480 228124 4 analog_io[26]
port 18 nsew signal bidirectional
rlabel metal3 s -960 175796 480 176036 4 analog_io[27]
port 19 nsew signal bidirectional
rlabel metal3 s -960 123572 480 123812 4 analog_io[28]
port 20 nsew signal bidirectional
rlabel metal3 s 583520 391628 584960 391868 6 analog_io[2]
port 21 nsew signal bidirectional
rlabel metal3 s 583520 444668 584960 444908 6 analog_io[3]
port 22 nsew signal bidirectional
rlabel metal3 s 583520 497844 584960 498084 6 analog_io[4]
port 23 nsew signal bidirectional
rlabel metal3 s 583520 551020 584960 551260 6 analog_io[5]
port 24 nsew signal bidirectional
rlabel metal3 s 583520 604060 584960 604300 6 analog_io[6]
port 25 nsew signal bidirectional
rlabel metal3 s 583520 657236 584960 657476 6 analog_io[7]
port 26 nsew signal bidirectional
rlabel metal2 s 575818 703520 575930 704960 6 analog_io[8]
port 27 nsew signal bidirectional
rlabel metal2 s 510958 703520 511070 704960 6 analog_io[9]
port 28 nsew signal bidirectional
rlabel metal3 s 583520 6476 584960 6716 6 io_in[0]
port 29 nsew signal input
rlabel metal3 s 583520 457996 584960 458236 6 io_in[10]
port 30 nsew signal input
rlabel metal3 s 583520 511172 584960 511412 6 io_in[11]
port 31 nsew signal input
rlabel metal3 s 583520 564212 584960 564452 6 io_in[12]
port 32 nsew signal input
rlabel metal3 s 583520 617388 584960 617628 6 io_in[13]
port 33 nsew signal input
rlabel metal3 s 583520 670564 584960 670804 6 io_in[14]
port 34 nsew signal input
rlabel metal2 s 559626 703520 559738 704960 6 io_in[15]
port 35 nsew signal input
rlabel metal2 s 494766 703520 494878 704960 6 io_in[16]
port 36 nsew signal input
rlabel metal2 s 429814 703520 429926 704960 6 io_in[17]
port 37 nsew signal input
rlabel metal2 s 364954 703520 365066 704960 6 io_in[18]
port 38 nsew signal input
rlabel metal2 s 300094 703520 300206 704960 6 io_in[19]
port 39 nsew signal input
rlabel metal3 s 583520 46188 584960 46428 6 io_in[1]
port 40 nsew signal input
rlabel metal2 s 235142 703520 235254 704960 6 io_in[20]
port 41 nsew signal input
rlabel metal2 s 170282 703520 170394 704960 6 io_in[21]
port 42 nsew signal input
rlabel metal2 s 105422 703520 105534 704960 6 io_in[22]
port 43 nsew signal input
rlabel metal2 s 40470 703520 40582 704960 6 io_in[23]
port 44 nsew signal input
rlabel metal3 s -960 684164 480 684404 4 io_in[24]
port 45 nsew signal input
rlabel metal3 s -960 631940 480 632180 4 io_in[25]
port 46 nsew signal input
rlabel metal3 s -960 579852 480 580092 4 io_in[26]
port 47 nsew signal input
rlabel metal3 s -960 527764 480 528004 4 io_in[27]
port 48 nsew signal input
rlabel metal3 s -960 475540 480 475780 4 io_in[28]
port 49 nsew signal input
rlabel metal3 s -960 423452 480 423692 4 io_in[29]
port 50 nsew signal input
rlabel metal3 s 583520 86036 584960 86276 6 io_in[2]
port 51 nsew signal input
rlabel metal3 s -960 371228 480 371468 4 io_in[30]
port 52 nsew signal input
rlabel metal3 s -960 319140 480 319380 4 io_in[31]
port 53 nsew signal input
rlabel metal3 s -960 267052 480 267292 4 io_in[32]
port 54 nsew signal input
rlabel metal3 s -960 214828 480 215068 4 io_in[33]
port 55 nsew signal input
rlabel metal3 s -960 162740 480 162980 4 io_in[34]
port 56 nsew signal input
rlabel metal3 s -960 110516 480 110756 4 io_in[35]
port 57 nsew signal input
rlabel metal3 s -960 71484 480 71724 4 io_in[36]
port 58 nsew signal input
rlabel metal3 s -960 32316 480 32556 4 io_in[37]
port 59 nsew signal input
rlabel metal3 s 583520 125884 584960 126124 6 io_in[3]
port 60 nsew signal input
rlabel metal3 s 583520 165732 584960 165972 6 io_in[4]
port 61 nsew signal input
rlabel metal3 s 583520 205580 584960 205820 6 io_in[5]
port 62 nsew signal input
rlabel metal3 s 583520 245428 584960 245668 6 io_in[6]
port 63 nsew signal input
rlabel metal3 s 583520 298604 584960 298844 6 io_in[7]
port 64 nsew signal input
rlabel metal3 s 583520 351780 584960 352020 6 io_in[8]
port 65 nsew signal input
rlabel metal3 s 583520 404820 584960 405060 6 io_in[9]
port 66 nsew signal input
rlabel metal3 s 583520 32996 584960 33236 6 io_oeb[0]
port 67 nsew signal tristate
rlabel metal3 s 583520 484516 584960 484756 6 io_oeb[10]
port 68 nsew signal tristate
rlabel metal3 s 583520 537692 584960 537932 6 io_oeb[11]
port 69 nsew signal tristate
rlabel metal3 s 583520 590868 584960 591108 6 io_oeb[12]
port 70 nsew signal tristate
rlabel metal3 s 583520 643908 584960 644148 6 io_oeb[13]
port 71 nsew signal tristate
rlabel metal3 s 583520 697084 584960 697324 6 io_oeb[14]
port 72 nsew signal tristate
rlabel metal2 s 527150 703520 527262 704960 6 io_oeb[15]
port 73 nsew signal tristate
rlabel metal2 s 462290 703520 462402 704960 6 io_oeb[16]
port 74 nsew signal tristate
rlabel metal2 s 397430 703520 397542 704960 6 io_oeb[17]
port 75 nsew signal tristate
rlabel metal2 s 332478 703520 332590 704960 6 io_oeb[18]
port 76 nsew signal tristate
rlabel metal2 s 267618 703520 267730 704960 6 io_oeb[19]
port 77 nsew signal tristate
rlabel metal3 s 583520 72844 584960 73084 6 io_oeb[1]
port 78 nsew signal tristate
rlabel metal2 s 202758 703520 202870 704960 6 io_oeb[20]
port 79 nsew signal tristate
rlabel metal2 s 137806 703520 137918 704960 6 io_oeb[21]
port 80 nsew signal tristate
rlabel metal2 s 72946 703520 73058 704960 6 io_oeb[22]
port 81 nsew signal tristate
rlabel metal2 s 8086 703520 8198 704960 6 io_oeb[23]
port 82 nsew signal tristate
rlabel metal3 s -960 658052 480 658292 4 io_oeb[24]
port 83 nsew signal tristate
rlabel metal3 s -960 605964 480 606204 4 io_oeb[25]
port 84 nsew signal tristate
rlabel metal3 s -960 553740 480 553980 4 io_oeb[26]
port 85 nsew signal tristate
rlabel metal3 s -960 501652 480 501892 4 io_oeb[27]
port 86 nsew signal tristate
rlabel metal3 s -960 449428 480 449668 4 io_oeb[28]
port 87 nsew signal tristate
rlabel metal3 s -960 397340 480 397580 4 io_oeb[29]
port 88 nsew signal tristate
rlabel metal3 s 583520 112692 584960 112932 6 io_oeb[2]
port 89 nsew signal tristate
rlabel metal3 s -960 345252 480 345492 4 io_oeb[30]
port 90 nsew signal tristate
rlabel metal3 s -960 293028 480 293268 4 io_oeb[31]
port 91 nsew signal tristate
rlabel metal3 s -960 240940 480 241180 4 io_oeb[32]
port 92 nsew signal tristate
rlabel metal3 s -960 188716 480 188956 4 io_oeb[33]
port 93 nsew signal tristate
rlabel metal3 s -960 136628 480 136868 4 io_oeb[34]
port 94 nsew signal tristate
rlabel metal3 s -960 84540 480 84780 4 io_oeb[35]
port 95 nsew signal tristate
rlabel metal3 s -960 45372 480 45612 4 io_oeb[36]
port 96 nsew signal tristate
rlabel metal3 s -960 6340 480 6580 4 io_oeb[37]
port 97 nsew signal tristate
rlabel metal3 s 583520 152540 584960 152780 6 io_oeb[3]
port 98 nsew signal tristate
rlabel metal3 s 583520 192388 584960 192628 6 io_oeb[4]
port 99 nsew signal tristate
rlabel metal3 s 583520 232236 584960 232476 6 io_oeb[5]
port 100 nsew signal tristate
rlabel metal3 s 583520 272084 584960 272324 6 io_oeb[6]
port 101 nsew signal tristate
rlabel metal3 s 583520 325124 584960 325364 6 io_oeb[7]
port 102 nsew signal tristate
rlabel metal3 s 583520 378300 584960 378540 6 io_oeb[8]
port 103 nsew signal tristate
rlabel metal3 s 583520 431476 584960 431716 6 io_oeb[9]
port 104 nsew signal tristate
rlabel metal3 s 583520 19668 584960 19908 6 io_out[0]
port 105 nsew signal tristate
rlabel metal3 s 583520 471324 584960 471564 6 io_out[10]
port 106 nsew signal tristate
rlabel metal3 s 583520 524364 584960 524604 6 io_out[11]
port 107 nsew signal tristate
rlabel metal3 s 583520 577540 584960 577780 6 io_out[12]
port 108 nsew signal tristate
rlabel metal3 s 583520 630716 584960 630956 6 io_out[13]
port 109 nsew signal tristate
rlabel metal3 s 583520 683756 584960 683996 6 io_out[14]
port 110 nsew signal tristate
rlabel metal2 s 543434 703520 543546 704960 6 io_out[15]
port 111 nsew signal tristate
rlabel metal2 s 478482 703520 478594 704960 6 io_out[16]
port 112 nsew signal tristate
rlabel metal2 s 413622 703520 413734 704960 6 io_out[17]
port 113 nsew signal tristate
rlabel metal2 s 348762 703520 348874 704960 6 io_out[18]
port 114 nsew signal tristate
rlabel metal2 s 283810 703520 283922 704960 6 io_out[19]
port 115 nsew signal tristate
rlabel metal3 s 583520 59516 584960 59756 6 io_out[1]
port 116 nsew signal tristate
rlabel metal2 s 218950 703520 219062 704960 6 io_out[20]
port 117 nsew signal tristate
rlabel metal2 s 154090 703520 154202 704960 6 io_out[21]
port 118 nsew signal tristate
rlabel metal2 s 89138 703520 89250 704960 6 io_out[22]
port 119 nsew signal tristate
rlabel metal2 s 24278 703520 24390 704960 6 io_out[23]
port 120 nsew signal tristate
rlabel metal3 s -960 671108 480 671348 4 io_out[24]
port 121 nsew signal tristate
rlabel metal3 s -960 619020 480 619260 4 io_out[25]
port 122 nsew signal tristate
rlabel metal3 s -960 566796 480 567036 4 io_out[26]
port 123 nsew signal tristate
rlabel metal3 s -960 514708 480 514948 4 io_out[27]
port 124 nsew signal tristate
rlabel metal3 s -960 462484 480 462724 4 io_out[28]
port 125 nsew signal tristate
rlabel metal3 s -960 410396 480 410636 4 io_out[29]
port 126 nsew signal tristate
rlabel metal3 s 583520 99364 584960 99604 6 io_out[2]
port 127 nsew signal tristate
rlabel metal3 s -960 358308 480 358548 4 io_out[30]
port 128 nsew signal tristate
rlabel metal3 s -960 306084 480 306324 4 io_out[31]
port 129 nsew signal tristate
rlabel metal3 s -960 253996 480 254236 4 io_out[32]
port 130 nsew signal tristate
rlabel metal3 s -960 201772 480 202012 4 io_out[33]
port 131 nsew signal tristate
rlabel metal3 s -960 149684 480 149924 4 io_out[34]
port 132 nsew signal tristate
rlabel metal3 s -960 97460 480 97700 4 io_out[35]
port 133 nsew signal tristate
rlabel metal3 s -960 58428 480 58668 4 io_out[36]
port 134 nsew signal tristate
rlabel metal3 s -960 19260 480 19500 4 io_out[37]
port 135 nsew signal tristate
rlabel metal3 s 583520 139212 584960 139452 6 io_out[3]
port 136 nsew signal tristate
rlabel metal3 s 583520 179060 584960 179300 6 io_out[4]
port 137 nsew signal tristate
rlabel metal3 s 583520 218908 584960 219148 6 io_out[5]
port 138 nsew signal tristate
rlabel metal3 s 583520 258756 584960 258996 6 io_out[6]
port 139 nsew signal tristate
rlabel metal3 s 583520 311932 584960 312172 6 io_out[7]
port 140 nsew signal tristate
rlabel metal3 s 583520 364972 584960 365212 6 io_out[8]
port 141 nsew signal tristate
rlabel metal3 s 583520 418148 584960 418388 6 io_out[9]
port 142 nsew signal tristate
rlabel metal2 s 125846 -960 125958 480 8 la_data_in[0]
port 143 nsew signal input
rlabel metal2 s 480506 -960 480618 480 8 la_data_in[100]
port 144 nsew signal input
rlabel metal2 s 484002 -960 484114 480 8 la_data_in[101]
port 145 nsew signal input
rlabel metal2 s 487590 -960 487702 480 8 la_data_in[102]
port 146 nsew signal input
rlabel metal2 s 491086 -960 491198 480 8 la_data_in[103]
port 147 nsew signal input
rlabel metal2 s 494674 -960 494786 480 8 la_data_in[104]
port 148 nsew signal input
rlabel metal2 s 498170 -960 498282 480 8 la_data_in[105]
port 149 nsew signal input
rlabel metal2 s 501758 -960 501870 480 8 la_data_in[106]
port 150 nsew signal input
rlabel metal2 s 505346 -960 505458 480 8 la_data_in[107]
port 151 nsew signal input
rlabel metal2 s 508842 -960 508954 480 8 la_data_in[108]
port 152 nsew signal input
rlabel metal2 s 512430 -960 512542 480 8 la_data_in[109]
port 153 nsew signal input
rlabel metal2 s 161266 -960 161378 480 8 la_data_in[10]
port 154 nsew signal input
rlabel metal2 s 515926 -960 516038 480 8 la_data_in[110]
port 155 nsew signal input
rlabel metal2 s 519514 -960 519626 480 8 la_data_in[111]
port 156 nsew signal input
rlabel metal2 s 523010 -960 523122 480 8 la_data_in[112]
port 157 nsew signal input
rlabel metal2 s 526598 -960 526710 480 8 la_data_in[113]
port 158 nsew signal input
rlabel metal2 s 530094 -960 530206 480 8 la_data_in[114]
port 159 nsew signal input
rlabel metal2 s 533682 -960 533794 480 8 la_data_in[115]
port 160 nsew signal input
rlabel metal2 s 537178 -960 537290 480 8 la_data_in[116]
port 161 nsew signal input
rlabel metal2 s 540766 -960 540878 480 8 la_data_in[117]
port 162 nsew signal input
rlabel metal2 s 544354 -960 544466 480 8 la_data_in[118]
port 163 nsew signal input
rlabel metal2 s 547850 -960 547962 480 8 la_data_in[119]
port 164 nsew signal input
rlabel metal2 s 164854 -960 164966 480 8 la_data_in[11]
port 165 nsew signal input
rlabel metal2 s 551438 -960 551550 480 8 la_data_in[120]
port 166 nsew signal input
rlabel metal2 s 554934 -960 555046 480 8 la_data_in[121]
port 167 nsew signal input
rlabel metal2 s 558522 -960 558634 480 8 la_data_in[122]
port 168 nsew signal input
rlabel metal2 s 562018 -960 562130 480 8 la_data_in[123]
port 169 nsew signal input
rlabel metal2 s 565606 -960 565718 480 8 la_data_in[124]
port 170 nsew signal input
rlabel metal2 s 569102 -960 569214 480 8 la_data_in[125]
port 171 nsew signal input
rlabel metal2 s 572690 -960 572802 480 8 la_data_in[126]
port 172 nsew signal input
rlabel metal2 s 576278 -960 576390 480 8 la_data_in[127]
port 173 nsew signal input
rlabel metal2 s 168350 -960 168462 480 8 la_data_in[12]
port 174 nsew signal input
rlabel metal2 s 171938 -960 172050 480 8 la_data_in[13]
port 175 nsew signal input
rlabel metal2 s 175434 -960 175546 480 8 la_data_in[14]
port 176 nsew signal input
rlabel metal2 s 179022 -960 179134 480 8 la_data_in[15]
port 177 nsew signal input
rlabel metal2 s 182518 -960 182630 480 8 la_data_in[16]
port 178 nsew signal input
rlabel metal2 s 186106 -960 186218 480 8 la_data_in[17]
port 179 nsew signal input
rlabel metal2 s 189694 -960 189806 480 8 la_data_in[18]
port 180 nsew signal input
rlabel metal2 s 193190 -960 193302 480 8 la_data_in[19]
port 181 nsew signal input
rlabel metal2 s 129342 -960 129454 480 8 la_data_in[1]
port 182 nsew signal input
rlabel metal2 s 196778 -960 196890 480 8 la_data_in[20]
port 183 nsew signal input
rlabel metal2 s 200274 -960 200386 480 8 la_data_in[21]
port 184 nsew signal input
rlabel metal2 s 203862 -960 203974 480 8 la_data_in[22]
port 185 nsew signal input
rlabel metal2 s 207358 -960 207470 480 8 la_data_in[23]
port 186 nsew signal input
rlabel metal2 s 210946 -960 211058 480 8 la_data_in[24]
port 187 nsew signal input
rlabel metal2 s 214442 -960 214554 480 8 la_data_in[25]
port 188 nsew signal input
rlabel metal2 s 218030 -960 218142 480 8 la_data_in[26]
port 189 nsew signal input
rlabel metal2 s 221526 -960 221638 480 8 la_data_in[27]
port 190 nsew signal input
rlabel metal2 s 225114 -960 225226 480 8 la_data_in[28]
port 191 nsew signal input
rlabel metal2 s 228702 -960 228814 480 8 la_data_in[29]
port 192 nsew signal input
rlabel metal2 s 132930 -960 133042 480 8 la_data_in[2]
port 193 nsew signal input
rlabel metal2 s 232198 -960 232310 480 8 la_data_in[30]
port 194 nsew signal input
rlabel metal2 s 235786 -960 235898 480 8 la_data_in[31]
port 195 nsew signal input
rlabel metal2 s 239282 -960 239394 480 8 la_data_in[32]
port 196 nsew signal input
rlabel metal2 s 242870 -960 242982 480 8 la_data_in[33]
port 197 nsew signal input
rlabel metal2 s 246366 -960 246478 480 8 la_data_in[34]
port 198 nsew signal input
rlabel metal2 s 249954 -960 250066 480 8 la_data_in[35]
port 199 nsew signal input
rlabel metal2 s 253450 -960 253562 480 8 la_data_in[36]
port 200 nsew signal input
rlabel metal2 s 257038 -960 257150 480 8 la_data_in[37]
port 201 nsew signal input
rlabel metal2 s 260626 -960 260738 480 8 la_data_in[38]
port 202 nsew signal input
rlabel metal2 s 264122 -960 264234 480 8 la_data_in[39]
port 203 nsew signal input
rlabel metal2 s 136426 -960 136538 480 8 la_data_in[3]
port 204 nsew signal input
rlabel metal2 s 267710 -960 267822 480 8 la_data_in[40]
port 205 nsew signal input
rlabel metal2 s 271206 -960 271318 480 8 la_data_in[41]
port 206 nsew signal input
rlabel metal2 s 274794 -960 274906 480 8 la_data_in[42]
port 207 nsew signal input
rlabel metal2 s 278290 -960 278402 480 8 la_data_in[43]
port 208 nsew signal input
rlabel metal2 s 281878 -960 281990 480 8 la_data_in[44]
port 209 nsew signal input
rlabel metal2 s 285374 -960 285486 480 8 la_data_in[45]
port 210 nsew signal input
rlabel metal2 s 288962 -960 289074 480 8 la_data_in[46]
port 211 nsew signal input
rlabel metal2 s 292550 -960 292662 480 8 la_data_in[47]
port 212 nsew signal input
rlabel metal2 s 296046 -960 296158 480 8 la_data_in[48]
port 213 nsew signal input
rlabel metal2 s 299634 -960 299746 480 8 la_data_in[49]
port 214 nsew signal input
rlabel metal2 s 140014 -960 140126 480 8 la_data_in[4]
port 215 nsew signal input
rlabel metal2 s 303130 -960 303242 480 8 la_data_in[50]
port 216 nsew signal input
rlabel metal2 s 306718 -960 306830 480 8 la_data_in[51]
port 217 nsew signal input
rlabel metal2 s 310214 -960 310326 480 8 la_data_in[52]
port 218 nsew signal input
rlabel metal2 s 313802 -960 313914 480 8 la_data_in[53]
port 219 nsew signal input
rlabel metal2 s 317298 -960 317410 480 8 la_data_in[54]
port 220 nsew signal input
rlabel metal2 s 320886 -960 320998 480 8 la_data_in[55]
port 221 nsew signal input
rlabel metal2 s 324382 -960 324494 480 8 la_data_in[56]
port 222 nsew signal input
rlabel metal2 s 327970 -960 328082 480 8 la_data_in[57]
port 223 nsew signal input
rlabel metal2 s 331558 -960 331670 480 8 la_data_in[58]
port 224 nsew signal input
rlabel metal2 s 335054 -960 335166 480 8 la_data_in[59]
port 225 nsew signal input
rlabel metal2 s 143510 -960 143622 480 8 la_data_in[5]
port 226 nsew signal input
rlabel metal2 s 338642 -960 338754 480 8 la_data_in[60]
port 227 nsew signal input
rlabel metal2 s 342138 -960 342250 480 8 la_data_in[61]
port 228 nsew signal input
rlabel metal2 s 345726 -960 345838 480 8 la_data_in[62]
port 229 nsew signal input
rlabel metal2 s 349222 -960 349334 480 8 la_data_in[63]
port 230 nsew signal input
rlabel metal2 s 352810 -960 352922 480 8 la_data_in[64]
port 231 nsew signal input
rlabel metal2 s 356306 -960 356418 480 8 la_data_in[65]
port 232 nsew signal input
rlabel metal2 s 359894 -960 360006 480 8 la_data_in[66]
port 233 nsew signal input
rlabel metal2 s 363482 -960 363594 480 8 la_data_in[67]
port 234 nsew signal input
rlabel metal2 s 366978 -960 367090 480 8 la_data_in[68]
port 235 nsew signal input
rlabel metal2 s 370566 -960 370678 480 8 la_data_in[69]
port 236 nsew signal input
rlabel metal2 s 147098 -960 147210 480 8 la_data_in[6]
port 237 nsew signal input
rlabel metal2 s 374062 -960 374174 480 8 la_data_in[70]
port 238 nsew signal input
rlabel metal2 s 377650 -960 377762 480 8 la_data_in[71]
port 239 nsew signal input
rlabel metal2 s 381146 -960 381258 480 8 la_data_in[72]
port 240 nsew signal input
rlabel metal2 s 384734 -960 384846 480 8 la_data_in[73]
port 241 nsew signal input
rlabel metal2 s 388230 -960 388342 480 8 la_data_in[74]
port 242 nsew signal input
rlabel metal2 s 391818 -960 391930 480 8 la_data_in[75]
port 243 nsew signal input
rlabel metal2 s 395314 -960 395426 480 8 la_data_in[76]
port 244 nsew signal input
rlabel metal2 s 398902 -960 399014 480 8 la_data_in[77]
port 245 nsew signal input
rlabel metal2 s 402490 -960 402602 480 8 la_data_in[78]
port 246 nsew signal input
rlabel metal2 s 405986 -960 406098 480 8 la_data_in[79]
port 247 nsew signal input
rlabel metal2 s 150594 -960 150706 480 8 la_data_in[7]
port 248 nsew signal input
rlabel metal2 s 409574 -960 409686 480 8 la_data_in[80]
port 249 nsew signal input
rlabel metal2 s 413070 -960 413182 480 8 la_data_in[81]
port 250 nsew signal input
rlabel metal2 s 416658 -960 416770 480 8 la_data_in[82]
port 251 nsew signal input
rlabel metal2 s 420154 -960 420266 480 8 la_data_in[83]
port 252 nsew signal input
rlabel metal2 s 423742 -960 423854 480 8 la_data_in[84]
port 253 nsew signal input
rlabel metal2 s 427238 -960 427350 480 8 la_data_in[85]
port 254 nsew signal input
rlabel metal2 s 430826 -960 430938 480 8 la_data_in[86]
port 255 nsew signal input
rlabel metal2 s 434414 -960 434526 480 8 la_data_in[87]
port 256 nsew signal input
rlabel metal2 s 437910 -960 438022 480 8 la_data_in[88]
port 257 nsew signal input
rlabel metal2 s 441498 -960 441610 480 8 la_data_in[89]
port 258 nsew signal input
rlabel metal2 s 154182 -960 154294 480 8 la_data_in[8]
port 259 nsew signal input
rlabel metal2 s 444994 -960 445106 480 8 la_data_in[90]
port 260 nsew signal input
rlabel metal2 s 448582 -960 448694 480 8 la_data_in[91]
port 261 nsew signal input
rlabel metal2 s 452078 -960 452190 480 8 la_data_in[92]
port 262 nsew signal input
rlabel metal2 s 455666 -960 455778 480 8 la_data_in[93]
port 263 nsew signal input
rlabel metal2 s 459162 -960 459274 480 8 la_data_in[94]
port 264 nsew signal input
rlabel metal2 s 462750 -960 462862 480 8 la_data_in[95]
port 265 nsew signal input
rlabel metal2 s 466246 -960 466358 480 8 la_data_in[96]
port 266 nsew signal input
rlabel metal2 s 469834 -960 469946 480 8 la_data_in[97]
port 267 nsew signal input
rlabel metal2 s 473422 -960 473534 480 8 la_data_in[98]
port 268 nsew signal input
rlabel metal2 s 476918 -960 477030 480 8 la_data_in[99]
port 269 nsew signal input
rlabel metal2 s 157770 -960 157882 480 8 la_data_in[9]
port 270 nsew signal input
rlabel metal2 s 126950 -960 127062 480 8 la_data_out[0]
port 271 nsew signal tristate
rlabel metal2 s 481702 -960 481814 480 8 la_data_out[100]
port 272 nsew signal tristate
rlabel metal2 s 485198 -960 485310 480 8 la_data_out[101]
port 273 nsew signal tristate
rlabel metal2 s 488786 -960 488898 480 8 la_data_out[102]
port 274 nsew signal tristate
rlabel metal2 s 492282 -960 492394 480 8 la_data_out[103]
port 275 nsew signal tristate
rlabel metal2 s 495870 -960 495982 480 8 la_data_out[104]
port 276 nsew signal tristate
rlabel metal2 s 499366 -960 499478 480 8 la_data_out[105]
port 277 nsew signal tristate
rlabel metal2 s 502954 -960 503066 480 8 la_data_out[106]
port 278 nsew signal tristate
rlabel metal2 s 506450 -960 506562 480 8 la_data_out[107]
port 279 nsew signal tristate
rlabel metal2 s 510038 -960 510150 480 8 la_data_out[108]
port 280 nsew signal tristate
rlabel metal2 s 513534 -960 513646 480 8 la_data_out[109]
port 281 nsew signal tristate
rlabel metal2 s 162462 -960 162574 480 8 la_data_out[10]
port 282 nsew signal tristate
rlabel metal2 s 517122 -960 517234 480 8 la_data_out[110]
port 283 nsew signal tristate
rlabel metal2 s 520710 -960 520822 480 8 la_data_out[111]
port 284 nsew signal tristate
rlabel metal2 s 524206 -960 524318 480 8 la_data_out[112]
port 285 nsew signal tristate
rlabel metal2 s 527794 -960 527906 480 8 la_data_out[113]
port 286 nsew signal tristate
rlabel metal2 s 531290 -960 531402 480 8 la_data_out[114]
port 287 nsew signal tristate
rlabel metal2 s 534878 -960 534990 480 8 la_data_out[115]
port 288 nsew signal tristate
rlabel metal2 s 538374 -960 538486 480 8 la_data_out[116]
port 289 nsew signal tristate
rlabel metal2 s 541962 -960 542074 480 8 la_data_out[117]
port 290 nsew signal tristate
rlabel metal2 s 545458 -960 545570 480 8 la_data_out[118]
port 291 nsew signal tristate
rlabel metal2 s 549046 -960 549158 480 8 la_data_out[119]
port 292 nsew signal tristate
rlabel metal2 s 166050 -960 166162 480 8 la_data_out[11]
port 293 nsew signal tristate
rlabel metal2 s 552634 -960 552746 480 8 la_data_out[120]
port 294 nsew signal tristate
rlabel metal2 s 556130 -960 556242 480 8 la_data_out[121]
port 295 nsew signal tristate
rlabel metal2 s 559718 -960 559830 480 8 la_data_out[122]
port 296 nsew signal tristate
rlabel metal2 s 563214 -960 563326 480 8 la_data_out[123]
port 297 nsew signal tristate
rlabel metal2 s 566802 -960 566914 480 8 la_data_out[124]
port 298 nsew signal tristate
rlabel metal2 s 570298 -960 570410 480 8 la_data_out[125]
port 299 nsew signal tristate
rlabel metal2 s 573886 -960 573998 480 8 la_data_out[126]
port 300 nsew signal tristate
rlabel metal2 s 577382 -960 577494 480 8 la_data_out[127]
port 301 nsew signal tristate
rlabel metal2 s 169546 -960 169658 480 8 la_data_out[12]
port 302 nsew signal tristate
rlabel metal2 s 173134 -960 173246 480 8 la_data_out[13]
port 303 nsew signal tristate
rlabel metal2 s 176630 -960 176742 480 8 la_data_out[14]
port 304 nsew signal tristate
rlabel metal2 s 180218 -960 180330 480 8 la_data_out[15]
port 305 nsew signal tristate
rlabel metal2 s 183714 -960 183826 480 8 la_data_out[16]
port 306 nsew signal tristate
rlabel metal2 s 187302 -960 187414 480 8 la_data_out[17]
port 307 nsew signal tristate
rlabel metal2 s 190798 -960 190910 480 8 la_data_out[18]
port 308 nsew signal tristate
rlabel metal2 s 194386 -960 194498 480 8 la_data_out[19]
port 309 nsew signal tristate
rlabel metal2 s 130538 -960 130650 480 8 la_data_out[1]
port 310 nsew signal tristate
rlabel metal2 s 197882 -960 197994 480 8 la_data_out[20]
port 311 nsew signal tristate
rlabel metal2 s 201470 -960 201582 480 8 la_data_out[21]
port 312 nsew signal tristate
rlabel metal2 s 205058 -960 205170 480 8 la_data_out[22]
port 313 nsew signal tristate
rlabel metal2 s 208554 -960 208666 480 8 la_data_out[23]
port 314 nsew signal tristate
rlabel metal2 s 212142 -960 212254 480 8 la_data_out[24]
port 315 nsew signal tristate
rlabel metal2 s 215638 -960 215750 480 8 la_data_out[25]
port 316 nsew signal tristate
rlabel metal2 s 219226 -960 219338 480 8 la_data_out[26]
port 317 nsew signal tristate
rlabel metal2 s 222722 -960 222834 480 8 la_data_out[27]
port 318 nsew signal tristate
rlabel metal2 s 226310 -960 226422 480 8 la_data_out[28]
port 319 nsew signal tristate
rlabel metal2 s 229806 -960 229918 480 8 la_data_out[29]
port 320 nsew signal tristate
rlabel metal2 s 134126 -960 134238 480 8 la_data_out[2]
port 321 nsew signal tristate
rlabel metal2 s 233394 -960 233506 480 8 la_data_out[30]
port 322 nsew signal tristate
rlabel metal2 s 236982 -960 237094 480 8 la_data_out[31]
port 323 nsew signal tristate
rlabel metal2 s 240478 -960 240590 480 8 la_data_out[32]
port 324 nsew signal tristate
rlabel metal2 s 244066 -960 244178 480 8 la_data_out[33]
port 325 nsew signal tristate
rlabel metal2 s 247562 -960 247674 480 8 la_data_out[34]
port 326 nsew signal tristate
rlabel metal2 s 251150 -960 251262 480 8 la_data_out[35]
port 327 nsew signal tristate
rlabel metal2 s 254646 -960 254758 480 8 la_data_out[36]
port 328 nsew signal tristate
rlabel metal2 s 258234 -960 258346 480 8 la_data_out[37]
port 329 nsew signal tristate
rlabel metal2 s 261730 -960 261842 480 8 la_data_out[38]
port 330 nsew signal tristate
rlabel metal2 s 265318 -960 265430 480 8 la_data_out[39]
port 331 nsew signal tristate
rlabel metal2 s 137622 -960 137734 480 8 la_data_out[3]
port 332 nsew signal tristate
rlabel metal2 s 268814 -960 268926 480 8 la_data_out[40]
port 333 nsew signal tristate
rlabel metal2 s 272402 -960 272514 480 8 la_data_out[41]
port 334 nsew signal tristate
rlabel metal2 s 275990 -960 276102 480 8 la_data_out[42]
port 335 nsew signal tristate
rlabel metal2 s 279486 -960 279598 480 8 la_data_out[43]
port 336 nsew signal tristate
rlabel metal2 s 283074 -960 283186 480 8 la_data_out[44]
port 337 nsew signal tristate
rlabel metal2 s 286570 -960 286682 480 8 la_data_out[45]
port 338 nsew signal tristate
rlabel metal2 s 290158 -960 290270 480 8 la_data_out[46]
port 339 nsew signal tristate
rlabel metal2 s 293654 -960 293766 480 8 la_data_out[47]
port 340 nsew signal tristate
rlabel metal2 s 297242 -960 297354 480 8 la_data_out[48]
port 341 nsew signal tristate
rlabel metal2 s 300738 -960 300850 480 8 la_data_out[49]
port 342 nsew signal tristate
rlabel metal2 s 141210 -960 141322 480 8 la_data_out[4]
port 343 nsew signal tristate
rlabel metal2 s 304326 -960 304438 480 8 la_data_out[50]
port 344 nsew signal tristate
rlabel metal2 s 307914 -960 308026 480 8 la_data_out[51]
port 345 nsew signal tristate
rlabel metal2 s 311410 -960 311522 480 8 la_data_out[52]
port 346 nsew signal tristate
rlabel metal2 s 314998 -960 315110 480 8 la_data_out[53]
port 347 nsew signal tristate
rlabel metal2 s 318494 -960 318606 480 8 la_data_out[54]
port 348 nsew signal tristate
rlabel metal2 s 322082 -960 322194 480 8 la_data_out[55]
port 349 nsew signal tristate
rlabel metal2 s 325578 -960 325690 480 8 la_data_out[56]
port 350 nsew signal tristate
rlabel metal2 s 329166 -960 329278 480 8 la_data_out[57]
port 351 nsew signal tristate
rlabel metal2 s 332662 -960 332774 480 8 la_data_out[58]
port 352 nsew signal tristate
rlabel metal2 s 336250 -960 336362 480 8 la_data_out[59]
port 353 nsew signal tristate
rlabel metal2 s 144706 -960 144818 480 8 la_data_out[5]
port 354 nsew signal tristate
rlabel metal2 s 339838 -960 339950 480 8 la_data_out[60]
port 355 nsew signal tristate
rlabel metal2 s 343334 -960 343446 480 8 la_data_out[61]
port 356 nsew signal tristate
rlabel metal2 s 346922 -960 347034 480 8 la_data_out[62]
port 357 nsew signal tristate
rlabel metal2 s 350418 -960 350530 480 8 la_data_out[63]
port 358 nsew signal tristate
rlabel metal2 s 354006 -960 354118 480 8 la_data_out[64]
port 359 nsew signal tristate
rlabel metal2 s 357502 -960 357614 480 8 la_data_out[65]
port 360 nsew signal tristate
rlabel metal2 s 361090 -960 361202 480 8 la_data_out[66]
port 361 nsew signal tristate
rlabel metal2 s 364586 -960 364698 480 8 la_data_out[67]
port 362 nsew signal tristate
rlabel metal2 s 368174 -960 368286 480 8 la_data_out[68]
port 363 nsew signal tristate
rlabel metal2 s 371670 -960 371782 480 8 la_data_out[69]
port 364 nsew signal tristate
rlabel metal2 s 148294 -960 148406 480 8 la_data_out[6]
port 365 nsew signal tristate
rlabel metal2 s 375258 -960 375370 480 8 la_data_out[70]
port 366 nsew signal tristate
rlabel metal2 s 378846 -960 378958 480 8 la_data_out[71]
port 367 nsew signal tristate
rlabel metal2 s 382342 -960 382454 480 8 la_data_out[72]
port 368 nsew signal tristate
rlabel metal2 s 385930 -960 386042 480 8 la_data_out[73]
port 369 nsew signal tristate
rlabel metal2 s 389426 -960 389538 480 8 la_data_out[74]
port 370 nsew signal tristate
rlabel metal2 s 393014 -960 393126 480 8 la_data_out[75]
port 371 nsew signal tristate
rlabel metal2 s 396510 -960 396622 480 8 la_data_out[76]
port 372 nsew signal tristate
rlabel metal2 s 400098 -960 400210 480 8 la_data_out[77]
port 373 nsew signal tristate
rlabel metal2 s 403594 -960 403706 480 8 la_data_out[78]
port 374 nsew signal tristate
rlabel metal2 s 407182 -960 407294 480 8 la_data_out[79]
port 375 nsew signal tristate
rlabel metal2 s 151790 -960 151902 480 8 la_data_out[7]
port 376 nsew signal tristate
rlabel metal2 s 410770 -960 410882 480 8 la_data_out[80]
port 377 nsew signal tristate
rlabel metal2 s 414266 -960 414378 480 8 la_data_out[81]
port 378 nsew signal tristate
rlabel metal2 s 417854 -960 417966 480 8 la_data_out[82]
port 379 nsew signal tristate
rlabel metal2 s 421350 -960 421462 480 8 la_data_out[83]
port 380 nsew signal tristate
rlabel metal2 s 424938 -960 425050 480 8 la_data_out[84]
port 381 nsew signal tristate
rlabel metal2 s 428434 -960 428546 480 8 la_data_out[85]
port 382 nsew signal tristate
rlabel metal2 s 432022 -960 432134 480 8 la_data_out[86]
port 383 nsew signal tristate
rlabel metal2 s 435518 -960 435630 480 8 la_data_out[87]
port 384 nsew signal tristate
rlabel metal2 s 439106 -960 439218 480 8 la_data_out[88]
port 385 nsew signal tristate
rlabel metal2 s 442602 -960 442714 480 8 la_data_out[89]
port 386 nsew signal tristate
rlabel metal2 s 155378 -960 155490 480 8 la_data_out[8]
port 387 nsew signal tristate
rlabel metal2 s 446190 -960 446302 480 8 la_data_out[90]
port 388 nsew signal tristate
rlabel metal2 s 449778 -960 449890 480 8 la_data_out[91]
port 389 nsew signal tristate
rlabel metal2 s 453274 -960 453386 480 8 la_data_out[92]
port 390 nsew signal tristate
rlabel metal2 s 456862 -960 456974 480 8 la_data_out[93]
port 391 nsew signal tristate
rlabel metal2 s 460358 -960 460470 480 8 la_data_out[94]
port 392 nsew signal tristate
rlabel metal2 s 463946 -960 464058 480 8 la_data_out[95]
port 393 nsew signal tristate
rlabel metal2 s 467442 -960 467554 480 8 la_data_out[96]
port 394 nsew signal tristate
rlabel metal2 s 471030 -960 471142 480 8 la_data_out[97]
port 395 nsew signal tristate
rlabel metal2 s 474526 -960 474638 480 8 la_data_out[98]
port 396 nsew signal tristate
rlabel metal2 s 478114 -960 478226 480 8 la_data_out[99]
port 397 nsew signal tristate
rlabel metal2 s 158874 -960 158986 480 8 la_data_out[9]
port 398 nsew signal tristate
rlabel metal2 s 128146 -960 128258 480 8 la_oenb[0]
port 399 nsew signal input
rlabel metal2 s 482806 -960 482918 480 8 la_oenb[100]
port 400 nsew signal input
rlabel metal2 s 486394 -960 486506 480 8 la_oenb[101]
port 401 nsew signal input
rlabel metal2 s 489890 -960 490002 480 8 la_oenb[102]
port 402 nsew signal input
rlabel metal2 s 493478 -960 493590 480 8 la_oenb[103]
port 403 nsew signal input
rlabel metal2 s 497066 -960 497178 480 8 la_oenb[104]
port 404 nsew signal input
rlabel metal2 s 500562 -960 500674 480 8 la_oenb[105]
port 405 nsew signal input
rlabel metal2 s 504150 -960 504262 480 8 la_oenb[106]
port 406 nsew signal input
rlabel metal2 s 507646 -960 507758 480 8 la_oenb[107]
port 407 nsew signal input
rlabel metal2 s 511234 -960 511346 480 8 la_oenb[108]
port 408 nsew signal input
rlabel metal2 s 514730 -960 514842 480 8 la_oenb[109]
port 409 nsew signal input
rlabel metal2 s 163658 -960 163770 480 8 la_oenb[10]
port 410 nsew signal input
rlabel metal2 s 518318 -960 518430 480 8 la_oenb[110]
port 411 nsew signal input
rlabel metal2 s 521814 -960 521926 480 8 la_oenb[111]
port 412 nsew signal input
rlabel metal2 s 525402 -960 525514 480 8 la_oenb[112]
port 413 nsew signal input
rlabel metal2 s 528990 -960 529102 480 8 la_oenb[113]
port 414 nsew signal input
rlabel metal2 s 532486 -960 532598 480 8 la_oenb[114]
port 415 nsew signal input
rlabel metal2 s 536074 -960 536186 480 8 la_oenb[115]
port 416 nsew signal input
rlabel metal2 s 539570 -960 539682 480 8 la_oenb[116]
port 417 nsew signal input
rlabel metal2 s 543158 -960 543270 480 8 la_oenb[117]
port 418 nsew signal input
rlabel metal2 s 546654 -960 546766 480 8 la_oenb[118]
port 419 nsew signal input
rlabel metal2 s 550242 -960 550354 480 8 la_oenb[119]
port 420 nsew signal input
rlabel metal2 s 167154 -960 167266 480 8 la_oenb[11]
port 421 nsew signal input
rlabel metal2 s 553738 -960 553850 480 8 la_oenb[120]
port 422 nsew signal input
rlabel metal2 s 557326 -960 557438 480 8 la_oenb[121]
port 423 nsew signal input
rlabel metal2 s 560822 -960 560934 480 8 la_oenb[122]
port 424 nsew signal input
rlabel metal2 s 564410 -960 564522 480 8 la_oenb[123]
port 425 nsew signal input
rlabel metal2 s 567998 -960 568110 480 8 la_oenb[124]
port 426 nsew signal input
rlabel metal2 s 571494 -960 571606 480 8 la_oenb[125]
port 427 nsew signal input
rlabel metal2 s 575082 -960 575194 480 8 la_oenb[126]
port 428 nsew signal input
rlabel metal2 s 578578 -960 578690 480 8 la_oenb[127]
port 429 nsew signal input
rlabel metal2 s 170742 -960 170854 480 8 la_oenb[12]
port 430 nsew signal input
rlabel metal2 s 174238 -960 174350 480 8 la_oenb[13]
port 431 nsew signal input
rlabel metal2 s 177826 -960 177938 480 8 la_oenb[14]
port 432 nsew signal input
rlabel metal2 s 181414 -960 181526 480 8 la_oenb[15]
port 433 nsew signal input
rlabel metal2 s 184910 -960 185022 480 8 la_oenb[16]
port 434 nsew signal input
rlabel metal2 s 188498 -960 188610 480 8 la_oenb[17]
port 435 nsew signal input
rlabel metal2 s 191994 -960 192106 480 8 la_oenb[18]
port 436 nsew signal input
rlabel metal2 s 195582 -960 195694 480 8 la_oenb[19]
port 437 nsew signal input
rlabel metal2 s 131734 -960 131846 480 8 la_oenb[1]
port 438 nsew signal input
rlabel metal2 s 199078 -960 199190 480 8 la_oenb[20]
port 439 nsew signal input
rlabel metal2 s 202666 -960 202778 480 8 la_oenb[21]
port 440 nsew signal input
rlabel metal2 s 206162 -960 206274 480 8 la_oenb[22]
port 441 nsew signal input
rlabel metal2 s 209750 -960 209862 480 8 la_oenb[23]
port 442 nsew signal input
rlabel metal2 s 213338 -960 213450 480 8 la_oenb[24]
port 443 nsew signal input
rlabel metal2 s 216834 -960 216946 480 8 la_oenb[25]
port 444 nsew signal input
rlabel metal2 s 220422 -960 220534 480 8 la_oenb[26]
port 445 nsew signal input
rlabel metal2 s 223918 -960 224030 480 8 la_oenb[27]
port 446 nsew signal input
rlabel metal2 s 227506 -960 227618 480 8 la_oenb[28]
port 447 nsew signal input
rlabel metal2 s 231002 -960 231114 480 8 la_oenb[29]
port 448 nsew signal input
rlabel metal2 s 135230 -960 135342 480 8 la_oenb[2]
port 449 nsew signal input
rlabel metal2 s 234590 -960 234702 480 8 la_oenb[30]
port 450 nsew signal input
rlabel metal2 s 238086 -960 238198 480 8 la_oenb[31]
port 451 nsew signal input
rlabel metal2 s 241674 -960 241786 480 8 la_oenb[32]
port 452 nsew signal input
rlabel metal2 s 245170 -960 245282 480 8 la_oenb[33]
port 453 nsew signal input
rlabel metal2 s 248758 -960 248870 480 8 la_oenb[34]
port 454 nsew signal input
rlabel metal2 s 252346 -960 252458 480 8 la_oenb[35]
port 455 nsew signal input
rlabel metal2 s 255842 -960 255954 480 8 la_oenb[36]
port 456 nsew signal input
rlabel metal2 s 259430 -960 259542 480 8 la_oenb[37]
port 457 nsew signal input
rlabel metal2 s 262926 -960 263038 480 8 la_oenb[38]
port 458 nsew signal input
rlabel metal2 s 266514 -960 266626 480 8 la_oenb[39]
port 459 nsew signal input
rlabel metal2 s 138818 -960 138930 480 8 la_oenb[3]
port 460 nsew signal input
rlabel metal2 s 270010 -960 270122 480 8 la_oenb[40]
port 461 nsew signal input
rlabel metal2 s 273598 -960 273710 480 8 la_oenb[41]
port 462 nsew signal input
rlabel metal2 s 277094 -960 277206 480 8 la_oenb[42]
port 463 nsew signal input
rlabel metal2 s 280682 -960 280794 480 8 la_oenb[43]
port 464 nsew signal input
rlabel metal2 s 284270 -960 284382 480 8 la_oenb[44]
port 465 nsew signal input
rlabel metal2 s 287766 -960 287878 480 8 la_oenb[45]
port 466 nsew signal input
rlabel metal2 s 291354 -960 291466 480 8 la_oenb[46]
port 467 nsew signal input
rlabel metal2 s 294850 -960 294962 480 8 la_oenb[47]
port 468 nsew signal input
rlabel metal2 s 298438 -960 298550 480 8 la_oenb[48]
port 469 nsew signal input
rlabel metal2 s 301934 -960 302046 480 8 la_oenb[49]
port 470 nsew signal input
rlabel metal2 s 142406 -960 142518 480 8 la_oenb[4]
port 471 nsew signal input
rlabel metal2 s 305522 -960 305634 480 8 la_oenb[50]
port 472 nsew signal input
rlabel metal2 s 309018 -960 309130 480 8 la_oenb[51]
port 473 nsew signal input
rlabel metal2 s 312606 -960 312718 480 8 la_oenb[52]
port 474 nsew signal input
rlabel metal2 s 316194 -960 316306 480 8 la_oenb[53]
port 475 nsew signal input
rlabel metal2 s 319690 -960 319802 480 8 la_oenb[54]
port 476 nsew signal input
rlabel metal2 s 323278 -960 323390 480 8 la_oenb[55]
port 477 nsew signal input
rlabel metal2 s 326774 -960 326886 480 8 la_oenb[56]
port 478 nsew signal input
rlabel metal2 s 330362 -960 330474 480 8 la_oenb[57]
port 479 nsew signal input
rlabel metal2 s 333858 -960 333970 480 8 la_oenb[58]
port 480 nsew signal input
rlabel metal2 s 337446 -960 337558 480 8 la_oenb[59]
port 481 nsew signal input
rlabel metal2 s 145902 -960 146014 480 8 la_oenb[5]
port 482 nsew signal input
rlabel metal2 s 340942 -960 341054 480 8 la_oenb[60]
port 483 nsew signal input
rlabel metal2 s 344530 -960 344642 480 8 la_oenb[61]
port 484 nsew signal input
rlabel metal2 s 348026 -960 348138 480 8 la_oenb[62]
port 485 nsew signal input
rlabel metal2 s 351614 -960 351726 480 8 la_oenb[63]
port 486 nsew signal input
rlabel metal2 s 355202 -960 355314 480 8 la_oenb[64]
port 487 nsew signal input
rlabel metal2 s 358698 -960 358810 480 8 la_oenb[65]
port 488 nsew signal input
rlabel metal2 s 362286 -960 362398 480 8 la_oenb[66]
port 489 nsew signal input
rlabel metal2 s 365782 -960 365894 480 8 la_oenb[67]
port 490 nsew signal input
rlabel metal2 s 369370 -960 369482 480 8 la_oenb[68]
port 491 nsew signal input
rlabel metal2 s 372866 -960 372978 480 8 la_oenb[69]
port 492 nsew signal input
rlabel metal2 s 149490 -960 149602 480 8 la_oenb[6]
port 493 nsew signal input
rlabel metal2 s 376454 -960 376566 480 8 la_oenb[70]
port 494 nsew signal input
rlabel metal2 s 379950 -960 380062 480 8 la_oenb[71]
port 495 nsew signal input
rlabel metal2 s 383538 -960 383650 480 8 la_oenb[72]
port 496 nsew signal input
rlabel metal2 s 387126 -960 387238 480 8 la_oenb[73]
port 497 nsew signal input
rlabel metal2 s 390622 -960 390734 480 8 la_oenb[74]
port 498 nsew signal input
rlabel metal2 s 394210 -960 394322 480 8 la_oenb[75]
port 499 nsew signal input
rlabel metal2 s 397706 -960 397818 480 8 la_oenb[76]
port 500 nsew signal input
rlabel metal2 s 401294 -960 401406 480 8 la_oenb[77]
port 501 nsew signal input
rlabel metal2 s 404790 -960 404902 480 8 la_oenb[78]
port 502 nsew signal input
rlabel metal2 s 408378 -960 408490 480 8 la_oenb[79]
port 503 nsew signal input
rlabel metal2 s 152986 -960 153098 480 8 la_oenb[7]
port 504 nsew signal input
rlabel metal2 s 411874 -960 411986 480 8 la_oenb[80]
port 505 nsew signal input
rlabel metal2 s 415462 -960 415574 480 8 la_oenb[81]
port 506 nsew signal input
rlabel metal2 s 418958 -960 419070 480 8 la_oenb[82]
port 507 nsew signal input
rlabel metal2 s 422546 -960 422658 480 8 la_oenb[83]
port 508 nsew signal input
rlabel metal2 s 426134 -960 426246 480 8 la_oenb[84]
port 509 nsew signal input
rlabel metal2 s 429630 -960 429742 480 8 la_oenb[85]
port 510 nsew signal input
rlabel metal2 s 433218 -960 433330 480 8 la_oenb[86]
port 511 nsew signal input
rlabel metal2 s 436714 -960 436826 480 8 la_oenb[87]
port 512 nsew signal input
rlabel metal2 s 440302 -960 440414 480 8 la_oenb[88]
port 513 nsew signal input
rlabel metal2 s 443798 -960 443910 480 8 la_oenb[89]
port 514 nsew signal input
rlabel metal2 s 156574 -960 156686 480 8 la_oenb[8]
port 515 nsew signal input
rlabel metal2 s 447386 -960 447498 480 8 la_oenb[90]
port 516 nsew signal input
rlabel metal2 s 450882 -960 450994 480 8 la_oenb[91]
port 517 nsew signal input
rlabel metal2 s 454470 -960 454582 480 8 la_oenb[92]
port 518 nsew signal input
rlabel metal2 s 458058 -960 458170 480 8 la_oenb[93]
port 519 nsew signal input
rlabel metal2 s 461554 -960 461666 480 8 la_oenb[94]
port 520 nsew signal input
rlabel metal2 s 465142 -960 465254 480 8 la_oenb[95]
port 521 nsew signal input
rlabel metal2 s 468638 -960 468750 480 8 la_oenb[96]
port 522 nsew signal input
rlabel metal2 s 472226 -960 472338 480 8 la_oenb[97]
port 523 nsew signal input
rlabel metal2 s 475722 -960 475834 480 8 la_oenb[98]
port 524 nsew signal input
rlabel metal2 s 479310 -960 479422 480 8 la_oenb[99]
port 525 nsew signal input
rlabel metal2 s 160070 -960 160182 480 8 la_oenb[9]
port 526 nsew signal input
rlabel metal2 s 579774 -960 579886 480 8 user_clock2
port 527 nsew signal input
rlabel metal2 s 580970 -960 581082 480 8 user_irq[0]
port 528 nsew signal tristate
rlabel metal2 s 582166 -960 582278 480 8 user_irq[1]
port 529 nsew signal tristate
rlabel metal2 s 583362 -960 583474 480 8 user_irq[2]
port 530 nsew signal tristate
rlabel metal5 s -2006 -934 585930 -314 8 vccd1
port 531 nsew power input
rlabel metal5 s -2966 2866 586890 3486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 38866 586890 39486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 74866 586890 75486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 110866 586890 111486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 146866 586890 147486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 182866 586890 183486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 218866 586890 219486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 254866 586890 255486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 290866 586890 291486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 326866 586890 327486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 362866 586890 363486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 398866 586890 399486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 434866 586890 435486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 470866 586890 471486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 506866 586890 507486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 542866 586890 543486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 578866 586890 579486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 614866 586890 615486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 650866 586890 651486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 686866 586890 687486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2006 704250 585930 704870 6 vccd1
port 531 nsew power input
rlabel metal4 s 181794 -1894 182414 198800 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 -1894 218414 198800 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 -1894 254414 198800 6 vccd1
port 531 nsew power input
rlabel metal4 s 289794 -1894 290414 198800 6 vccd1
port 531 nsew power input
rlabel metal4 s 325794 -1894 326414 198800 6 vccd1
port 531 nsew power input
rlabel metal4 s 361794 -1894 362414 198800 6 vccd1
port 531 nsew power input
rlabel metal4 s 397794 -1894 398414 198800 6 vccd1
port 531 nsew power input
rlabel metal4 s -2006 -934 -1386 704870 4 vccd1
port 531 nsew power input
rlabel metal4 s 585310 -934 585930 704870 6 vccd1
port 531 nsew power input
rlabel metal4 s 1794 -1894 2414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 37794 -1894 38414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 -1894 74414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 -1894 110414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 -1894 146414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 181794 509939 182414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 509939 218414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 509939 254414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 289794 509939 290414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 325794 509939 326414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 361794 509939 362414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 397794 509939 398414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 433794 -1894 434414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 469794 -1894 470414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 505794 -1894 506414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 541794 -1894 542414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 577794 -1894 578414 705830 6 vccd1
port 531 nsew power input
rlabel metal5 s -3926 -2854 587850 -2234 8 vccd2
port 532 nsew power input
rlabel metal5 s -4886 6586 588810 7206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 42586 588810 43206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 78586 588810 79206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 114586 588810 115206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 150586 588810 151206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 186586 588810 187206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 222586 588810 223206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 258586 588810 259206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 294586 588810 295206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 330586 588810 331206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 366586 588810 367206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 402586 588810 403206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 438586 588810 439206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 474586 588810 475206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 510586 588810 511206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 546586 588810 547206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 582586 588810 583206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 618586 588810 619206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 654586 588810 655206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 690586 588810 691206 6 vccd2
port 532 nsew power input
rlabel metal5 s -3926 706170 587850 706790 6 vccd2
port 532 nsew power input
rlabel metal4 s 185514 -3814 186134 198800 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 -3814 222134 198800 6 vccd2
port 532 nsew power input
rlabel metal4 s 257514 -3814 258134 198800 6 vccd2
port 532 nsew power input
rlabel metal4 s 293514 -3814 294134 198800 6 vccd2
port 532 nsew power input
rlabel metal4 s 329514 -3814 330134 198800 6 vccd2
port 532 nsew power input
rlabel metal4 s 365514 -3814 366134 198800 6 vccd2
port 532 nsew power input
rlabel metal4 s 401514 -3814 402134 198800 6 vccd2
port 532 nsew power input
rlabel metal4 s -3926 -2854 -3306 706790 4 vccd2
port 532 nsew power input
rlabel metal4 s 587230 -2854 587850 706790 6 vccd2
port 532 nsew power input
rlabel metal4 s 5514 -3814 6134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 41514 -3814 42134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 -3814 78134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 -3814 114134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 149514 -3814 150134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 185514 509939 186134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 509939 222134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 257514 509939 258134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 293514 509939 294134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 329514 509939 330134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 365514 509939 366134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 401514 509939 402134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 437514 -3814 438134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 473514 -3814 474134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 509514 -3814 510134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 545514 -3814 546134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 581514 -3814 582134 707750 6 vccd2
port 532 nsew power input
rlabel metal5 s -5846 -4774 589770 -4154 8 vdda1
port 533 nsew power input
rlabel metal5 s -6806 10306 590730 10926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 46306 590730 46926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 82306 590730 82926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 118306 590730 118926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 154306 590730 154926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 190306 590730 190926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 226306 590730 226926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 262306 590730 262926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 298306 590730 298926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 334306 590730 334926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 370306 590730 370926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 406306 590730 406926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 442306 590730 442926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 478306 590730 478926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 514306 590730 514926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 550306 590730 550926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 586306 590730 586926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 622306 590730 622926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 658306 590730 658926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 694306 590730 694926 6 vdda1
port 533 nsew power input
rlabel metal5 s -5846 708090 589770 708710 6 vdda1
port 533 nsew power input
rlabel metal4 s 189234 -5734 189854 198800 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 -5734 225854 198800 6 vdda1
port 533 nsew power input
rlabel metal4 s 261234 -5734 261854 198800 6 vdda1
port 533 nsew power input
rlabel metal4 s 297234 -5734 297854 198800 6 vdda1
port 533 nsew power input
rlabel metal4 s 333234 -5734 333854 198800 6 vdda1
port 533 nsew power input
rlabel metal4 s 369234 -5734 369854 198800 6 vdda1
port 533 nsew power input
rlabel metal4 s 405234 -5734 405854 198800 6 vdda1
port 533 nsew power input
rlabel metal4 s -5846 -4774 -5226 708710 4 vdda1
port 533 nsew power input
rlabel metal4 s 589150 -4774 589770 708710 6 vdda1
port 533 nsew power input
rlabel metal4 s 9234 -5734 9854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 45234 -5734 45854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 -5734 81854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 -5734 117854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 153234 -5734 153854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 189234 509939 189854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 509939 225854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 261234 509939 261854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 297234 509939 297854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 333234 509939 333854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 369234 509939 369854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 405234 509939 405854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 441234 -5734 441854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 477234 -5734 477854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 513234 -5734 513854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 549234 -5734 549854 709670 6 vdda1
port 533 nsew power input
rlabel metal5 s -7766 -6694 591690 -6074 8 vdda2
port 534 nsew power input
rlabel metal5 s -8726 14026 592650 14646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 50026 592650 50646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 86026 592650 86646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 122026 592650 122646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 158026 592650 158646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 194026 592650 194646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 230026 592650 230646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 266026 592650 266646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 302026 592650 302646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 338026 592650 338646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 374026 592650 374646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 410026 592650 410646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 446026 592650 446646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 482026 592650 482646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 518026 592650 518646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 554026 592650 554646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 590026 592650 590646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 626026 592650 626646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 662026 592650 662646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 698026 592650 698646 6 vdda2
port 534 nsew power input
rlabel metal5 s -7766 710010 591690 710630 6 vdda2
port 534 nsew power input
rlabel metal4 s 192954 -7654 193574 198800 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 -7654 229574 198800 6 vdda2
port 534 nsew power input
rlabel metal4 s 264954 -7654 265574 198800 6 vdda2
port 534 nsew power input
rlabel metal4 s 300954 -7654 301574 198800 6 vdda2
port 534 nsew power input
rlabel metal4 s 336954 -7654 337574 198800 6 vdda2
port 534 nsew power input
rlabel metal4 s 372954 -7654 373574 198800 6 vdda2
port 534 nsew power input
rlabel metal4 s 408954 -7654 409574 198800 6 vdda2
port 534 nsew power input
rlabel metal4 s -7766 -6694 -7146 710630 4 vdda2
port 534 nsew power input
rlabel metal4 s 591070 -6694 591690 710630 6 vdda2
port 534 nsew power input
rlabel metal4 s 12954 -7654 13574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 48954 -7654 49574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 -7654 85574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 120954 -7654 121574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 156954 -7654 157574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 192954 509939 193574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 509939 229574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 264954 509939 265574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 300954 509939 301574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 336954 509939 337574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 372954 509939 373574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 408954 509939 409574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 444954 -7654 445574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 480954 -7654 481574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 516954 -7654 517574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 552954 -7654 553574 711590 6 vdda2
port 534 nsew power input
rlabel metal5 s -6806 -5734 590730 -5114 8 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 28306 590730 28926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 64306 590730 64926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 100306 590730 100926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 136306 590730 136926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 172306 590730 172926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 208306 590730 208926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 244306 590730 244926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 280306 590730 280926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 316306 590730 316926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 352306 590730 352926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 388306 590730 388926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 424306 590730 424926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 460306 590730 460926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 496306 590730 496926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 532306 590730 532926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 568306 590730 568926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 604306 590730 604926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 640306 590730 640926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 676306 590730 676926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 709050 590730 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 171234 -5734 171854 198800 6 vssa1
port 535 nsew ground input
rlabel metal4 s 207234 -5734 207854 198800 6 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 -5734 243854 198800 6 vssa1
port 535 nsew ground input
rlabel metal4 s 279234 -5734 279854 198800 6 vssa1
port 535 nsew ground input
rlabel metal4 s 315234 -5734 315854 198800 6 vssa1
port 535 nsew ground input
rlabel metal4 s 351234 -5734 351854 198800 6 vssa1
port 535 nsew ground input
rlabel metal4 s 387234 -5734 387854 198800 6 vssa1
port 535 nsew ground input
rlabel metal4 s -6806 -5734 -6186 709670 4 vssa1
port 535 nsew ground input
rlabel metal4 s 27234 -5734 27854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 63234 -5734 63854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 -5734 99854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 135234 -5734 135854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 171234 509939 171854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 207234 509939 207854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 509939 243854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 279234 509939 279854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 315234 509939 315854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 351234 509939 351854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 387234 509939 387854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 423234 -5734 423854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 459234 -5734 459854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 495234 -5734 495854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 531234 -5734 531854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 567234 -5734 567854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 590110 -5734 590730 709670 6 vssa1
port 535 nsew ground input
rlabel metal5 s -8726 -7654 592650 -7034 8 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 32026 592650 32646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 68026 592650 68646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 104026 592650 104646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 140026 592650 140646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 176026 592650 176646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 212026 592650 212646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 248026 592650 248646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 284026 592650 284646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 320026 592650 320646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 356026 592650 356646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 392026 592650 392646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 428026 592650 428646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 464026 592650 464646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 500026 592650 500646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 536026 592650 536646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 572026 592650 572646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 608026 592650 608646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 644026 592650 644646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 680026 592650 680646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 710970 592650 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 174954 -7654 175574 198800 6 vssa2
port 536 nsew ground input
rlabel metal4 s 210954 -7654 211574 198800 6 vssa2
port 536 nsew ground input
rlabel metal4 s 246954 -7654 247574 198800 6 vssa2
port 536 nsew ground input
rlabel metal4 s 282954 -7654 283574 198800 6 vssa2
port 536 nsew ground input
rlabel metal4 s 318954 -7654 319574 198800 6 vssa2
port 536 nsew ground input
rlabel metal4 s 354954 -7654 355574 198800 6 vssa2
port 536 nsew ground input
rlabel metal4 s 390954 -7654 391574 198800 6 vssa2
port 536 nsew ground input
rlabel metal4 s -8726 -7654 -8106 711590 4 vssa2
port 536 nsew ground input
rlabel metal4 s 30954 -7654 31574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 -7654 67574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 -7654 103574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 138954 -7654 139574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 174954 509939 175574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 210954 509939 211574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 246954 509939 247574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 282954 509939 283574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 318954 509939 319574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 354954 509939 355574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 390954 509939 391574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 426954 -7654 427574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 462954 -7654 463574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 498954 -7654 499574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 534954 -7654 535574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 570954 -7654 571574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 592030 -7654 592650 711590 6 vssa2
port 536 nsew ground input
rlabel metal5 s -2966 -1894 586890 -1274 8 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 20866 586890 21486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 56866 586890 57486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 92866 586890 93486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 128866 586890 129486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 164866 586890 165486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 200866 586890 201486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 236866 586890 237486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 272866 586890 273486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 308866 586890 309486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 344866 586890 345486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 380866 586890 381486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 416866 586890 417486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 452866 586890 453486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 488866 586890 489486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 524866 586890 525486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 560866 586890 561486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 596866 586890 597486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 632866 586890 633486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 668866 586890 669486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 705210 586890 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 163794 -1894 164414 198800 6 vssd1
port 537 nsew ground input
rlabel metal4 s 199794 -1894 200414 198800 6 vssd1
port 537 nsew ground input
rlabel metal4 s 235794 -1894 236414 198800 6 vssd1
port 537 nsew ground input
rlabel metal4 s 271794 -1894 272414 198800 6 vssd1
port 537 nsew ground input
rlabel metal4 s 307794 -1894 308414 198800 6 vssd1
port 537 nsew ground input
rlabel metal4 s 343794 -1894 344414 198800 6 vssd1
port 537 nsew ground input
rlabel metal4 s 379794 -1894 380414 198800 6 vssd1
port 537 nsew ground input
rlabel metal4 s 415794 -1894 416414 198800 6 vssd1
port 537 nsew ground input
rlabel metal4 s -2966 -1894 -2346 705830 4 vssd1
port 537 nsew ground input
rlabel metal4 s 19794 -1894 20414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 55794 -1894 56414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 -1894 92414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 127794 -1894 128414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 163794 509939 164414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 199794 509939 200414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 235794 509939 236414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 271794 509939 272414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 307794 509939 308414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 343794 509939 344414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 379794 509939 380414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 415794 509939 416414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 451794 -1894 452414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 487794 -1894 488414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 523794 -1894 524414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 559794 -1894 560414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 586270 -1894 586890 705830 6 vssd1
port 537 nsew ground input
rlabel metal5 s -4886 -3814 588810 -3194 8 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 24586 588810 25206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 60586 588810 61206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 96586 588810 97206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 132586 588810 133206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 168586 588810 169206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 204586 588810 205206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 240586 588810 241206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 276586 588810 277206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 312586 588810 313206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 348586 588810 349206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 384586 588810 385206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 420586 588810 421206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 456586 588810 457206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 492586 588810 493206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 528586 588810 529206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 564586 588810 565206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 600586 588810 601206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 636586 588810 637206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 672586 588810 673206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 707130 588810 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 167514 -3814 168134 198800 6 vssd2
port 538 nsew ground input
rlabel metal4 s 203514 -3814 204134 198800 6 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 -3814 240134 198800 6 vssd2
port 538 nsew ground input
rlabel metal4 s 275514 -3814 276134 198800 6 vssd2
port 538 nsew ground input
rlabel metal4 s 311514 -3814 312134 198800 6 vssd2
port 538 nsew ground input
rlabel metal4 s 347514 -3814 348134 198800 6 vssd2
port 538 nsew ground input
rlabel metal4 s 383514 -3814 384134 198800 6 vssd2
port 538 nsew ground input
rlabel metal4 s 419514 -3814 420134 198800 6 vssd2
port 538 nsew ground input
rlabel metal4 s -4886 -3814 -4266 707750 4 vssd2
port 538 nsew ground input
rlabel metal4 s 23514 -3814 24134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 59514 -3814 60134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 -3814 96134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 131514 -3814 132134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 167514 509939 168134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 203514 509939 204134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 509939 240134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 275514 509939 276134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 311514 509939 312134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 347514 509939 348134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 383514 509939 384134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 419514 509939 420134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 455514 -3814 456134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 491514 -3814 492134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 527514 -3814 528134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 563514 -3814 564134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 588190 -3814 588810 707750 6 vssd2
port 538 nsew ground input
rlabel metal2 s 542 -960 654 480 8 wb_clk_i
port 539 nsew signal input
rlabel metal2 s 1646 -960 1758 480 8 wb_rst_i
port 540 nsew signal input
rlabel metal2 s 2842 -960 2954 480 8 wbs_ack_o
port 541 nsew signal tristate
rlabel metal2 s 7626 -960 7738 480 8 wbs_adr_i[0]
port 542 nsew signal input
rlabel metal2 s 47830 -960 47942 480 8 wbs_adr_i[10]
port 543 nsew signal input
rlabel metal2 s 51326 -960 51438 480 8 wbs_adr_i[11]
port 544 nsew signal input
rlabel metal2 s 54914 -960 55026 480 8 wbs_adr_i[12]
port 545 nsew signal input
rlabel metal2 s 58410 -960 58522 480 8 wbs_adr_i[13]
port 546 nsew signal input
rlabel metal2 s 61998 -960 62110 480 8 wbs_adr_i[14]
port 547 nsew signal input
rlabel metal2 s 65494 -960 65606 480 8 wbs_adr_i[15]
port 548 nsew signal input
rlabel metal2 s 69082 -960 69194 480 8 wbs_adr_i[16]
port 549 nsew signal input
rlabel metal2 s 72578 -960 72690 480 8 wbs_adr_i[17]
port 550 nsew signal input
rlabel metal2 s 76166 -960 76278 480 8 wbs_adr_i[18]
port 551 nsew signal input
rlabel metal2 s 79662 -960 79774 480 8 wbs_adr_i[19]
port 552 nsew signal input
rlabel metal2 s 12318 -960 12430 480 8 wbs_adr_i[1]
port 553 nsew signal input
rlabel metal2 s 83250 -960 83362 480 8 wbs_adr_i[20]
port 554 nsew signal input
rlabel metal2 s 86838 -960 86950 480 8 wbs_adr_i[21]
port 555 nsew signal input
rlabel metal2 s 90334 -960 90446 480 8 wbs_adr_i[22]
port 556 nsew signal input
rlabel metal2 s 93922 -960 94034 480 8 wbs_adr_i[23]
port 557 nsew signal input
rlabel metal2 s 97418 -960 97530 480 8 wbs_adr_i[24]
port 558 nsew signal input
rlabel metal2 s 101006 -960 101118 480 8 wbs_adr_i[25]
port 559 nsew signal input
rlabel metal2 s 104502 -960 104614 480 8 wbs_adr_i[26]
port 560 nsew signal input
rlabel metal2 s 108090 -960 108202 480 8 wbs_adr_i[27]
port 561 nsew signal input
rlabel metal2 s 111586 -960 111698 480 8 wbs_adr_i[28]
port 562 nsew signal input
rlabel metal2 s 115174 -960 115286 480 8 wbs_adr_i[29]
port 563 nsew signal input
rlabel metal2 s 17010 -960 17122 480 8 wbs_adr_i[2]
port 564 nsew signal input
rlabel metal2 s 118762 -960 118874 480 8 wbs_adr_i[30]
port 565 nsew signal input
rlabel metal2 s 122258 -960 122370 480 8 wbs_adr_i[31]
port 566 nsew signal input
rlabel metal2 s 21794 -960 21906 480 8 wbs_adr_i[3]
port 567 nsew signal input
rlabel metal2 s 26486 -960 26598 480 8 wbs_adr_i[4]
port 568 nsew signal input
rlabel metal2 s 30074 -960 30186 480 8 wbs_adr_i[5]
port 569 nsew signal input
rlabel metal2 s 33570 -960 33682 480 8 wbs_adr_i[6]
port 570 nsew signal input
rlabel metal2 s 37158 -960 37270 480 8 wbs_adr_i[7]
port 571 nsew signal input
rlabel metal2 s 40654 -960 40766 480 8 wbs_adr_i[8]
port 572 nsew signal input
rlabel metal2 s 44242 -960 44354 480 8 wbs_adr_i[9]
port 573 nsew signal input
rlabel metal2 s 4038 -960 4150 480 8 wbs_cyc_i
port 574 nsew signal input
rlabel metal2 s 8730 -960 8842 480 8 wbs_dat_i[0]
port 575 nsew signal input
rlabel metal2 s 48934 -960 49046 480 8 wbs_dat_i[10]
port 576 nsew signal input
rlabel metal2 s 52522 -960 52634 480 8 wbs_dat_i[11]
port 577 nsew signal input
rlabel metal2 s 56018 -960 56130 480 8 wbs_dat_i[12]
port 578 nsew signal input
rlabel metal2 s 59606 -960 59718 480 8 wbs_dat_i[13]
port 579 nsew signal input
rlabel metal2 s 63194 -960 63306 480 8 wbs_dat_i[14]
port 580 nsew signal input
rlabel metal2 s 66690 -960 66802 480 8 wbs_dat_i[15]
port 581 nsew signal input
rlabel metal2 s 70278 -960 70390 480 8 wbs_dat_i[16]
port 582 nsew signal input
rlabel metal2 s 73774 -960 73886 480 8 wbs_dat_i[17]
port 583 nsew signal input
rlabel metal2 s 77362 -960 77474 480 8 wbs_dat_i[18]
port 584 nsew signal input
rlabel metal2 s 80858 -960 80970 480 8 wbs_dat_i[19]
port 585 nsew signal input
rlabel metal2 s 13514 -960 13626 480 8 wbs_dat_i[1]
port 586 nsew signal input
rlabel metal2 s 84446 -960 84558 480 8 wbs_dat_i[20]
port 587 nsew signal input
rlabel metal2 s 87942 -960 88054 480 8 wbs_dat_i[21]
port 588 nsew signal input
rlabel metal2 s 91530 -960 91642 480 8 wbs_dat_i[22]
port 589 nsew signal input
rlabel metal2 s 95118 -960 95230 480 8 wbs_dat_i[23]
port 590 nsew signal input
rlabel metal2 s 98614 -960 98726 480 8 wbs_dat_i[24]
port 591 nsew signal input
rlabel metal2 s 102202 -960 102314 480 8 wbs_dat_i[25]
port 592 nsew signal input
rlabel metal2 s 105698 -960 105810 480 8 wbs_dat_i[26]
port 593 nsew signal input
rlabel metal2 s 109286 -960 109398 480 8 wbs_dat_i[27]
port 594 nsew signal input
rlabel metal2 s 112782 -960 112894 480 8 wbs_dat_i[28]
port 595 nsew signal input
rlabel metal2 s 116370 -960 116482 480 8 wbs_dat_i[29]
port 596 nsew signal input
rlabel metal2 s 18206 -960 18318 480 8 wbs_dat_i[2]
port 597 nsew signal input
rlabel metal2 s 119866 -960 119978 480 8 wbs_dat_i[30]
port 598 nsew signal input
rlabel metal2 s 123454 -960 123566 480 8 wbs_dat_i[31]
port 599 nsew signal input
rlabel metal2 s 22990 -960 23102 480 8 wbs_dat_i[3]
port 600 nsew signal input
rlabel metal2 s 27682 -960 27794 480 8 wbs_dat_i[4]
port 601 nsew signal input
rlabel metal2 s 31270 -960 31382 480 8 wbs_dat_i[5]
port 602 nsew signal input
rlabel metal2 s 34766 -960 34878 480 8 wbs_dat_i[6]
port 603 nsew signal input
rlabel metal2 s 38354 -960 38466 480 8 wbs_dat_i[7]
port 604 nsew signal input
rlabel metal2 s 41850 -960 41962 480 8 wbs_dat_i[8]
port 605 nsew signal input
rlabel metal2 s 45438 -960 45550 480 8 wbs_dat_i[9]
port 606 nsew signal input
rlabel metal2 s 9926 -960 10038 480 8 wbs_dat_o[0]
port 607 nsew signal tristate
rlabel metal2 s 50130 -960 50242 480 8 wbs_dat_o[10]
port 608 nsew signal tristate
rlabel metal2 s 53718 -960 53830 480 8 wbs_dat_o[11]
port 609 nsew signal tristate
rlabel metal2 s 57214 -960 57326 480 8 wbs_dat_o[12]
port 610 nsew signal tristate
rlabel metal2 s 60802 -960 60914 480 8 wbs_dat_o[13]
port 611 nsew signal tristate
rlabel metal2 s 64298 -960 64410 480 8 wbs_dat_o[14]
port 612 nsew signal tristate
rlabel metal2 s 67886 -960 67998 480 8 wbs_dat_o[15]
port 613 nsew signal tristate
rlabel metal2 s 71474 -960 71586 480 8 wbs_dat_o[16]
port 614 nsew signal tristate
rlabel metal2 s 74970 -960 75082 480 8 wbs_dat_o[17]
port 615 nsew signal tristate
rlabel metal2 s 78558 -960 78670 480 8 wbs_dat_o[18]
port 616 nsew signal tristate
rlabel metal2 s 82054 -960 82166 480 8 wbs_dat_o[19]
port 617 nsew signal tristate
rlabel metal2 s 14710 -960 14822 480 8 wbs_dat_o[1]
port 618 nsew signal tristate
rlabel metal2 s 85642 -960 85754 480 8 wbs_dat_o[20]
port 619 nsew signal tristate
rlabel metal2 s 89138 -960 89250 480 8 wbs_dat_o[21]
port 620 nsew signal tristate
rlabel metal2 s 92726 -960 92838 480 8 wbs_dat_o[22]
port 621 nsew signal tristate
rlabel metal2 s 96222 -960 96334 480 8 wbs_dat_o[23]
port 622 nsew signal tristate
rlabel metal2 s 99810 -960 99922 480 8 wbs_dat_o[24]
port 623 nsew signal tristate
rlabel metal2 s 103306 -960 103418 480 8 wbs_dat_o[25]
port 624 nsew signal tristate
rlabel metal2 s 106894 -960 107006 480 8 wbs_dat_o[26]
port 625 nsew signal tristate
rlabel metal2 s 110482 -960 110594 480 8 wbs_dat_o[27]
port 626 nsew signal tristate
rlabel metal2 s 113978 -960 114090 480 8 wbs_dat_o[28]
port 627 nsew signal tristate
rlabel metal2 s 117566 -960 117678 480 8 wbs_dat_o[29]
port 628 nsew signal tristate
rlabel metal2 s 19402 -960 19514 480 8 wbs_dat_o[2]
port 629 nsew signal tristate
rlabel metal2 s 121062 -960 121174 480 8 wbs_dat_o[30]
port 630 nsew signal tristate
rlabel metal2 s 124650 -960 124762 480 8 wbs_dat_o[31]
port 631 nsew signal tristate
rlabel metal2 s 24186 -960 24298 480 8 wbs_dat_o[3]
port 632 nsew signal tristate
rlabel metal2 s 28878 -960 28990 480 8 wbs_dat_o[4]
port 633 nsew signal tristate
rlabel metal2 s 32374 -960 32486 480 8 wbs_dat_o[5]
port 634 nsew signal tristate
rlabel metal2 s 35962 -960 36074 480 8 wbs_dat_o[6]
port 635 nsew signal tristate
rlabel metal2 s 39550 -960 39662 480 8 wbs_dat_o[7]
port 636 nsew signal tristate
rlabel metal2 s 43046 -960 43158 480 8 wbs_dat_o[8]
port 637 nsew signal tristate
rlabel metal2 s 46634 -960 46746 480 8 wbs_dat_o[9]
port 638 nsew signal tristate
rlabel metal2 s 11122 -960 11234 480 8 wbs_sel_i[0]
port 639 nsew signal input
rlabel metal2 s 15906 -960 16018 480 8 wbs_sel_i[1]
port 640 nsew signal input
rlabel metal2 s 20598 -960 20710 480 8 wbs_sel_i[2]
port 641 nsew signal input
rlabel metal2 s 25290 -960 25402 480 8 wbs_sel_i[3]
port 642 nsew signal input
rlabel metal2 s 5234 -960 5346 480 8 wbs_stb_i
port 643 nsew signal input
rlabel metal2 s 6430 -960 6542 480 8 wbs_we_i
port 644 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
